module DivSqrtRawFN_small_e23_s489(
  input          clock,
  input          reset,
  output         io_inReady,
  input          io_inValid,
  input          io_a_isNaN,
  input          io_a_isInf,
  input          io_a_isZero,
  input          io_a_sign,
  input  [24:0]  io_a_sExp,
  input  [489:0] io_a_sig,
  input          io_b_isNaN,
  input          io_b_isInf,
  input          io_b_isZero,
  input          io_b_sign,
  input  [24:0]  io_b_sExp,
  input  [489:0] io_b_sig,
  input  [2:0]   io_roundingMode,
  output         io_rawOutValid_div,
  output [2:0]   io_roundingModeOut,
  output         io_invalidExc,
  output         io_infiniteExc,
  output         io_rawOut_isNaN,
  output         io_rawOut_isInf,
  output         io_rawOut_isZero,
  output         io_rawOut_sign,
  output [24:0]  io_rawOut_sExp,
  output [491:0] io_rawOut_sig
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [511:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [511:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] cycleNum; // @[DivSqrtRecFN_small.scala 224:33]
  reg  inReady; // @[DivSqrtRecFN_small.scala 225:33]
  reg  rawOutValid; // @[DivSqrtRecFN_small.scala 226:33]
  reg  majorExc_Z; // @[DivSqrtRecFN_small.scala 229:29]
  reg  isNaN_Z; // @[DivSqrtRecFN_small.scala 231:29]
  reg  isInf_Z; // @[DivSqrtRecFN_small.scala 232:29]
  reg  isZero_Z; // @[DivSqrtRecFN_small.scala 233:29]
  reg  sign_Z; // @[DivSqrtRecFN_small.scala 234:29]
  reg [24:0] sExp_Z; // @[DivSqrtRecFN_small.scala 235:29]
  reg [488:0] fractB_Z; // @[DivSqrtRecFN_small.scala 236:29]
  reg [2:0] roundingMode_Z; // @[DivSqrtRecFN_small.scala 237:29]
  reg [490:0] rem_Z; // @[DivSqrtRecFN_small.scala 243:29]
  reg  notZeroRem_Z; // @[DivSqrtRecFN_small.scala 244:29]
  reg [490:0] sigX_Z; // @[DivSqrtRecFN_small.scala 245:29]
  wire  notSigNaNIn_invalidExc_S_div = io_a_isZero & io_b_isZero | io_a_isInf & io_b_isInf; // @[DivSqrtRecFN_small.scala 254:42]
  wire  _notSigNaNIn_invalidExc_S_sqrt_T = ~io_a_isNaN; // @[DivSqrtRecFN_small.scala 256:9]
  wire  _majorExc_S_T_2 = io_a_isNaN & ~io_a_sig[487]; // @[common.scala 82:46]
  wire  _majorExc_S_T_9 = io_b_isNaN & ~io_b_sig[487]; // @[common.scala 82:46]
  wire  _majorExc_S_T_11 = _majorExc_S_T_2 | _majorExc_S_T_9 | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 260:66]
  wire  _majorExc_S_T_15 = _notSigNaNIn_invalidExc_S_sqrt_T & ~io_a_isInf & io_b_isZero; // @[DivSqrtRecFN_small.scala 262:51]
  wire  majorExc_S = _majorExc_S_T_11 | _majorExc_S_T_15; // @[DivSqrtRecFN_small.scala 261:46]
  wire  isNaN_S = io_a_isNaN | io_b_isNaN | notSigNaNIn_invalidExc_S_div; // @[DivSqrtRecFN_small.scala 267:42]
  wire  isInf_S = io_a_isInf | io_b_isZero; // @[DivSqrtRecFN_small.scala 269:63]
  wire  isZero_S = io_a_isZero | io_b_isInf; // @[DivSqrtRecFN_small.scala 270:64]
  wire  sign_S = io_a_sign ^ io_b_sign; // @[DivSqrtRecFN_small.scala 271:30]
  wire  specialCaseA_S = io_a_isNaN | io_a_isInf | io_a_isZero; // @[DivSqrtRecFN_small.scala 273:55]
  wire  specialCaseB_S = io_b_isNaN | io_b_isInf | io_b_isZero; // @[DivSqrtRecFN_small.scala 274:55]
  wire  normalCase_S_div = ~specialCaseA_S & ~specialCaseB_S; // @[DivSqrtRecFN_small.scala 275:45]
  wire [22:0] _sExpQuot_S_div_T_2 = ~io_b_sExp[22:0]; // @[DivSqrtRecFN_small.scala 281:40]
  wire [23:0] _sExpQuot_S_div_T_4 = {io_b_sExp[23],_sExpQuot_S_div_T_2}; // @[DivSqrtRecFN_small.scala 281:71]
  wire [24:0] _GEN_15 = {{1{_sExpQuot_S_div_T_4[23]}},_sExpQuot_S_div_T_4}; // @[DivSqrtRecFN_small.scala 280:21]
  wire [25:0] sExpQuot_S_div = $signed(io_a_sExp) + $signed(_GEN_15); // @[DivSqrtRecFN_small.scala 280:21]
  wire [3:0] _sSatExpQuot_S_div_T_2 = 26'she00000 <= $signed(sExpQuot_S_div) ? 4'h6 : sExpQuot_S_div[24:21]; // @[DivSqrtRecFN_small.scala 284:16]
  wire [24:0] sSatExpQuot_S_div = {_sSatExpQuot_S_div_T_2,sExpQuot_S_div[20:0]}; // @[DivSqrtRecFN_small.scala 289:11]
  wire  idle = cycleNum == 9'h0; // @[DivSqrtRecFN_small.scala 296:25]
  wire  entering = inReady & io_inValid; // @[DivSqrtRecFN_small.scala 297:28]
  wire  entering_normalCase = entering & normalCase_S_div; // @[DivSqrtRecFN_small.scala 298:40]
  wire  skipCycle2 = cycleNum == 9'h3 & sigX_Z[490]; // @[DivSqrtRecFN_small.scala 301:39]
  wire  _inReady_T_1 = entering & ~normalCase_S_div; // @[DivSqrtRecFN_small.scala 305:26]
  wire [8:0] _inReady_T_17 = cycleNum - 9'h1; // @[DivSqrtRecFN_small.scala 313:56]
  wire  _inReady_T_18 = _inReady_T_17 <= 9'h1; // @[DivSqrtRecFN_small.scala 317:38]
  wire  _inReady_T_19 = ~entering & ~skipCycle2 & _inReady_T_18; // @[DivSqrtRecFN_small.scala 313:16]
  wire  _inReady_T_20 = _inReady_T_1 | _inReady_T_19; // @[DivSqrtRecFN_small.scala 312:15]
  wire  _inReady_T_23 = _inReady_T_20 | skipCycle2; // @[DivSqrtRecFN_small.scala 313:95]
  wire  _rawOutValid_T_18 = _inReady_T_17 == 9'h1; // @[DivSqrtRecFN_small.scala 318:42]
  wire  _rawOutValid_T_19 = ~entering & ~skipCycle2 & _rawOutValid_T_18; // @[DivSqrtRecFN_small.scala 313:16]
  wire  _rawOutValid_T_20 = _inReady_T_1 | _rawOutValid_T_19; // @[DivSqrtRecFN_small.scala 312:15]
  wire  _rawOutValid_T_23 = _rawOutValid_T_20 | skipCycle2; // @[DivSqrtRecFN_small.scala 313:95]
  wire [8:0] _cycleNum_T_6 = entering_normalCase ? 9'h1eb : 9'h0; // @[DivSqrtRecFN_small.scala 306:16]
  wire [8:0] _GEN_16 = {{8'd0}, _inReady_T_1}; // @[DivSqrtRecFN_small.scala 305:57]
  wire [8:0] _cycleNum_T_7 = _GEN_16 | _cycleNum_T_6; // @[DivSqrtRecFN_small.scala 305:57]
  wire [8:0] _cycleNum_T_14 = ~entering & ~skipCycle2 ? _inReady_T_17 : 9'h0; // @[DivSqrtRecFN_small.scala 313:16]
  wire [8:0] _cycleNum_T_15 = _cycleNum_T_7 | _cycleNum_T_14; // @[DivSqrtRecFN_small.scala 312:15]
  wire [8:0] _GEN_17 = {{8'd0}, skipCycle2}; // @[DivSqrtRecFN_small.scala 313:95]
  wire [8:0] _cycleNum_T_17 = _cycleNum_T_15 | _GEN_17; // @[DivSqrtRecFN_small.scala 313:95]
  wire  _GEN_0 = ~idle | entering ? _inReady_T_23 : inReady; // @[DivSqrtRecFN_small.scala 303:31 317:17 225:33]
  wire  _T_2 = ~inReady; // @[DivSqrtRecFN_small.scala 340:23]
  wire [488:0] _fractB_Z_T_3 = {io_b_sig[487:0], 1'h0}; // @[DivSqrtRecFN_small.scala 342:90]
  wire [488:0] _fractB_Z_T_4 = inReady ? _fractB_Z_T_3 : 489'h0; // @[DivSqrtRecFN_small.scala 342:16]
  wire [487:0] _fractB_Z_T_25 = _T_2 ? fractB_Z[488:1] : 488'h0; // @[DivSqrtRecFN_small.scala 346:16]
  wire [488:0] _GEN_18 = {{1'd0}, _fractB_Z_T_25}; // @[DivSqrtRecFN_small.scala 345:100]
  wire [488:0] _fractB_Z_T_26 = _fractB_Z_T_4 | _GEN_18; // @[DivSqrtRecFN_small.scala 345:100]
  wire [490:0] _rem_T_2 = {io_a_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 352:47]
  wire [490:0] _rem_T_3 = inReady ? _rem_T_2 : 491'h0; // @[DivSqrtRecFN_small.scala 352:12]
  wire [491:0] _rem_T_12 = {{1'd0}, _rem_T_3}; // @[DivSqrtRecFN_small.scala 352:57]
  wire [491:0] _rem_T_14 = {rem_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 359:29]
  wire [491:0] _rem_T_15 = _T_2 ? _rem_T_14 : 492'h0; // @[DivSqrtRecFN_small.scala 359:12]
  wire [491:0] rem = _rem_T_12 | _rem_T_15; // @[DivSqrtRecFN_small.scala 358:11]
  wire [511:0] _bitMask_T = 512'h1 << cycleNum; // @[DivSqrtRecFN_small.scala 360:23]
  wire [509:0] bitMask = _bitMask_T[511:2]; // @[DivSqrtRecFN_small.scala 360:34]
  wire [490:0] _trialTerm_T_2 = {io_b_sig, 1'h0}; // @[DivSqrtRecFN_small.scala 362:48]
  wire [490:0] _trialTerm_T_3 = inReady ? _trialTerm_T_2 : 491'h0; // @[DivSqrtRecFN_small.scala 362:12]
  wire [488:0] _trialTerm_T_11 = _T_2 ? fractB_Z : 489'h0; // @[DivSqrtRecFN_small.scala 365:12]
  wire [490:0] _GEN_19 = {{2'd0}, _trialTerm_T_11}; // @[DivSqrtRecFN_small.scala 364:74]
  wire [490:0] _trialTerm_T_12 = _trialTerm_T_3 | _GEN_19; // @[DivSqrtRecFN_small.scala 364:74]
  wire [489:0] _trialTerm_T_17 = _T_2 ? 490'h200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
     : 490'h0; // @[DivSqrtRecFN_small.scala 366:12]
  wire [490:0] _GEN_20 = {{1'd0}, _trialTerm_T_17}; // @[DivSqrtRecFN_small.scala 365:74]
  wire [490:0] _trialTerm_T_18 = _trialTerm_T_12 | _GEN_20; // @[DivSqrtRecFN_small.scala 365:74]
  wire [491:0] _trialTerm_T_21 = {sigX_Z, 1'h0}; // @[DivSqrtRecFN_small.scala 367:44]
  wire [491:0] trialTerm = {{1'd0}, _trialTerm_T_18}; // @[DivSqrtRecFN_small.scala 366:74]
  wire [492:0] _trialRem_T = {1'b0,$signed(rem)}; // @[DivSqrtRecFN_small.scala 368:24]
  wire [492:0] _trialRem_T_1 = {1'b0,$signed(trialTerm)}; // @[DivSqrtRecFN_small.scala 368:42]
  wire [493:0] trialRem = $signed(_trialRem_T) - $signed(_trialRem_T_1); // @[DivSqrtRecFN_small.scala 368:29]
  wire  newBit = 494'sh0 <= $signed(trialRem); // @[DivSqrtRecFN_small.scala 369:23]
  wire [493:0] _nextRem_Z_T = $signed(_trialRem_T) - $signed(_trialRem_T_1); // @[DivSqrtRecFN_small.scala 371:42]
  wire [493:0] _nextRem_Z_T_1 = newBit ? _nextRem_Z_T : {{2'd0}, rem}; // @[DivSqrtRecFN_small.scala 371:24]
  wire [490:0] nextRem_Z = _nextRem_Z_T_1[490:0]; // @[DivSqrtRecFN_small.scala 371:54]
  wire [490:0] _sigX_Z_T_2 = {newBit, 490'h0}; // @[DivSqrtRecFN_small.scala 394:50]
  wire [490:0] _sigX_Z_T_3 = inReady ? _sigX_Z_T_2 : 491'h0; // @[DivSqrtRecFN_small.scala 394:16]
  wire [490:0] _sigX_Z_T_12 = _T_2 ? sigX_Z : 491'h0; // @[DivSqrtRecFN_small.scala 397:16]
  wire [490:0] _sigX_Z_T_13 = _sigX_Z_T_3 | _sigX_Z_T_12; // @[DivSqrtRecFN_small.scala 396:74]
  wire [509:0] _sigX_Z_T_16 = _T_2 & newBit ? bitMask : 510'h0; // @[DivSqrtRecFN_small.scala 398:16]
  wire [509:0] _GEN_25 = {{19'd0}, _sigX_Z_T_13}; // @[DivSqrtRecFN_small.scala 397:74]
  wire [509:0] _sigX_Z_T_17 = _GEN_25 | _sigX_Z_T_16; // @[DivSqrtRecFN_small.scala 397:74]
  wire [509:0] _GEN_14 = entering | _T_2 ? _sigX_Z_T_17 : {{19'd0}, sigX_Z}; // @[DivSqrtRecFN_small.scala 390:34 393:16 245:29]
  wire [491:0] _GEN_26 = {{491'd0}, notZeroRem_Z}; // @[DivSqrtRecFN_small.scala 414:35]
  assign io_inReady = inReady; // @[DivSqrtRecFN_small.scala 322:16]
  assign io_rawOutValid_div = rawOutValid; // @[DivSqrtRecFN_small.scala 404:40]
  assign io_roundingModeOut = roundingMode_Z; // @[DivSqrtRecFN_small.scala 406:25]
  assign io_invalidExc = majorExc_Z & isNaN_Z; // @[DivSqrtRecFN_small.scala 407:36]
  assign io_infiniteExc = majorExc_Z & ~isNaN_Z; // @[DivSqrtRecFN_small.scala 408:36]
  assign io_rawOut_isNaN = isNaN_Z; // @[DivSqrtRecFN_small.scala 409:22]
  assign io_rawOut_isInf = isInf_Z; // @[DivSqrtRecFN_small.scala 410:22]
  assign io_rawOut_isZero = isZero_Z; // @[DivSqrtRecFN_small.scala 411:22]
  assign io_rawOut_sign = sign_Z; // @[DivSqrtRecFN_small.scala 412:22]
  assign io_rawOut_sExp = sExp_Z; // @[DivSqrtRecFN_small.scala 413:22]
  assign io_rawOut_sig = _trialTerm_T_21 | _GEN_26; // @[DivSqrtRecFN_small.scala 414:35]
  always @(posedge clock) begin
    if (reset) begin // @[DivSqrtRecFN_small.scala 224:33]
      cycleNum <= 9'h0; // @[DivSqrtRecFN_small.scala 224:33]
    end else if (~idle | entering) begin // @[DivSqrtRecFN_small.scala 303:31]
      cycleNum <= _cycleNum_T_17; // @[DivSqrtRecFN_small.scala 319:18]
    end
    inReady <= reset | _GEN_0; // @[DivSqrtRecFN_small.scala 225:{33,33}]
    if (reset) begin // @[DivSqrtRecFN_small.scala 226:33]
      rawOutValid <= 1'h0; // @[DivSqrtRecFN_small.scala 226:33]
    end else if (~idle | entering) begin // @[DivSqrtRecFN_small.scala 303:31]
      rawOutValid <= _rawOutValid_T_23; // @[DivSqrtRecFN_small.scala 318:21]
    end
    if (entering) begin // @[DivSqrtRecFN_small.scala 326:21]
      majorExc_Z <= majorExc_S; // @[DivSqrtRecFN_small.scala 328:20]
    end
    if (entering) begin // @[DivSqrtRecFN_small.scala 326:21]
      isNaN_Z <= isNaN_S; // @[DivSqrtRecFN_small.scala 329:20]
    end
    if (entering) begin // @[DivSqrtRecFN_small.scala 326:21]
      isInf_Z <= isInf_S; // @[DivSqrtRecFN_small.scala 330:20]
    end
    if (entering) begin // @[DivSqrtRecFN_small.scala 326:21]
      isZero_Z <= isZero_S; // @[DivSqrtRecFN_small.scala 331:20]
    end
    if (entering) begin // @[DivSqrtRecFN_small.scala 326:21]
      sign_Z <= sign_S; // @[DivSqrtRecFN_small.scala 332:20]
    end
    if (entering) begin // @[DivSqrtRecFN_small.scala 326:21]
      sExp_Z <= sSatExpQuot_S_div; // @[DivSqrtRecFN_small.scala 333:16]
    end
    if (entering) begin // @[DivSqrtRecFN_small.scala 340:46]
      fractB_Z <= _fractB_Z_T_26; // @[DivSqrtRecFN_small.scala 341:18]
    end
    if (entering) begin // @[DivSqrtRecFN_small.scala 326:21]
      roundingMode_Z <= io_roundingMode; // @[DivSqrtRecFN_small.scala 338:24]
    end
    if (entering | _T_2) begin // @[DivSqrtRecFN_small.scala 390:34]
      rem_Z <= nextRem_Z; // @[DivSqrtRecFN_small.scala 392:15]
    end
    if (entering | _T_2) begin // @[DivSqrtRecFN_small.scala 390:34]
      if (inReady | newBit) begin // @[DivSqrtRecFN_small.scala 380:31]
        notZeroRem_Z <= $signed(trialRem) != 494'sh0;
      end
    end
    sigX_Z <= _GEN_14[490:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleNum = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  inReady = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rawOutValid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  majorExc_Z = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  isNaN_Z = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  isInf_Z = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  isZero_Z = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sign_Z = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sExp_Z = _RAND_8[24:0];
  _RAND_9 = {16{`RANDOM}};
  fractB_Z = _RAND_9[488:0];
  _RAND_10 = {1{`RANDOM}};
  roundingMode_Z = _RAND_10[2:0];
  _RAND_11 = {16{`RANDOM}};
  rem_Z = _RAND_11[490:0];
  _RAND_12 = {1{`RANDOM}};
  notZeroRem_Z = _RAND_12[0:0];
  _RAND_13 = {16{`RANDOM}};
  sigX_Z = _RAND_13[490:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DivSqrtRecFMToRaw_small_e23_s489(
  input          clock,
  input          reset,
  output         io_inReady,
  input          io_inValid,
  input  [512:0] io_a,
  input  [512:0] io_b,
  input  [2:0]   io_roundingMode,
  output         io_rawOutValid_div,
  output [2:0]   io_roundingModeOut,
  output         io_invalidExc,
  output         io_infiniteExc,
  output         io_rawOut_isNaN,
  output         io_rawOut_isInf,
  output         io_rawOut_isZero,
  output         io_rawOut_sign,
  output [24:0]  io_rawOut_sExp,
  output [491:0] io_rawOut_sig
);
  wire  divSqrtRawFN__clock; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__reset; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_inReady; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_inValid; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_a_isNaN; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_a_isInf; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_a_isZero; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_a_sign; // @[DivSqrtRecFN_small.scala 446:15]
  wire [24:0] divSqrtRawFN__io_a_sExp; // @[DivSqrtRecFN_small.scala 446:15]
  wire [489:0] divSqrtRawFN__io_a_sig; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_b_isNaN; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_b_isInf; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_b_isZero; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_b_sign; // @[DivSqrtRecFN_small.scala 446:15]
  wire [24:0] divSqrtRawFN__io_b_sExp; // @[DivSqrtRecFN_small.scala 446:15]
  wire [489:0] divSqrtRawFN__io_b_sig; // @[DivSqrtRecFN_small.scala 446:15]
  wire [2:0] divSqrtRawFN__io_roundingMode; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 446:15]
  wire [2:0] divSqrtRawFN__io_roundingModeOut; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_invalidExc; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_infiniteExc; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 446:15]
  wire  divSqrtRawFN__io_rawOut_sign; // @[DivSqrtRecFN_small.scala 446:15]
  wire [24:0] divSqrtRawFN__io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 446:15]
  wire [491:0] divSqrtRawFN__io_rawOut_sig; // @[DivSqrtRecFN_small.scala 446:15]
  wire [23:0] divSqrtRawFN_io_a_exp = io_a[511:488]; // @[rawFloatFromRecFN.scala 51:21]
  wire  divSqrtRawFN_io_a_isZero = divSqrtRawFN_io_a_exp[23:21] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  divSqrtRawFN_io_a_isSpecial = divSqrtRawFN_io_a_exp[23:22] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _divSqrtRawFN_io_a_out_sig_T = ~divSqrtRawFN_io_a_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _divSqrtRawFN_io_a_out_sig_T_1 = {1'h0,_divSqrtRawFN_io_a_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  wire [23:0] divSqrtRawFN_io_b_exp = io_b[511:488]; // @[rawFloatFromRecFN.scala 51:21]
  wire  divSqrtRawFN_io_b_isZero = divSqrtRawFN_io_b_exp[23:21] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  divSqrtRawFN_io_b_isSpecial = divSqrtRawFN_io_b_exp[23:22] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  _divSqrtRawFN_io_b_out_sig_T = ~divSqrtRawFN_io_b_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [1:0] _divSqrtRawFN_io_b_out_sig_T_1 = {1'h0,_divSqrtRawFN_io_b_out_sig_T}; // @[rawFloatFromRecFN.scala 61:32]
  DivSqrtRawFN_small_e23_s489 divSqrtRawFN_ ( // @[DivSqrtRecFN_small.scala 446:15]
    .clock(divSqrtRawFN__clock),
    .reset(divSqrtRawFN__reset),
    .io_inReady(divSqrtRawFN__io_inReady),
    .io_inValid(divSqrtRawFN__io_inValid),
    .io_a_isNaN(divSqrtRawFN__io_a_isNaN),
    .io_a_isInf(divSqrtRawFN__io_a_isInf),
    .io_a_isZero(divSqrtRawFN__io_a_isZero),
    .io_a_sign(divSqrtRawFN__io_a_sign),
    .io_a_sExp(divSqrtRawFN__io_a_sExp),
    .io_a_sig(divSqrtRawFN__io_a_sig),
    .io_b_isNaN(divSqrtRawFN__io_b_isNaN),
    .io_b_isInf(divSqrtRawFN__io_b_isInf),
    .io_b_isZero(divSqrtRawFN__io_b_isZero),
    .io_b_sign(divSqrtRawFN__io_b_sign),
    .io_b_sExp(divSqrtRawFN__io_b_sExp),
    .io_b_sig(divSqrtRawFN__io_b_sig),
    .io_roundingMode(divSqrtRawFN__io_roundingMode),
    .io_rawOutValid_div(divSqrtRawFN__io_rawOutValid_div),
    .io_roundingModeOut(divSqrtRawFN__io_roundingModeOut),
    .io_invalidExc(divSqrtRawFN__io_invalidExc),
    .io_infiniteExc(divSqrtRawFN__io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRawFN__io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRawFN__io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRawFN__io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRawFN__io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRawFN__io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRawFN__io_rawOut_sig)
  );
  assign io_inReady = divSqrtRawFN__io_inReady; // @[DivSqrtRecFN_small.scala 448:16]
  assign io_rawOutValid_div = divSqrtRawFN__io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 455:25]
  assign io_roundingModeOut = divSqrtRawFN__io_roundingModeOut; // @[DivSqrtRecFN_small.scala 457:25]
  assign io_invalidExc = divSqrtRawFN__io_invalidExc; // @[DivSqrtRecFN_small.scala 458:25]
  assign io_infiniteExc = divSqrtRawFN__io_infiniteExc; // @[DivSqrtRecFN_small.scala 459:25]
  assign io_rawOut_isNaN = divSqrtRawFN__io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 460:25]
  assign io_rawOut_isInf = divSqrtRawFN__io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 460:25]
  assign io_rawOut_isZero = divSqrtRawFN__io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 460:25]
  assign io_rawOut_sign = divSqrtRawFN__io_rawOut_sign; // @[DivSqrtRecFN_small.scala 460:25]
  assign io_rawOut_sExp = divSqrtRawFN__io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 460:25]
  assign io_rawOut_sig = divSqrtRawFN__io_rawOut_sig; // @[DivSqrtRecFN_small.scala 460:25]
  assign divSqrtRawFN__clock = clock;
  assign divSqrtRawFN__reset = reset;
  assign divSqrtRawFN__io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 449:34]
  assign divSqrtRawFN__io_a_isNaN = divSqrtRawFN_io_a_isSpecial & divSqrtRawFN_io_a_exp[21]; // @[rawFloatFromRecFN.scala 56:33]
  assign divSqrtRawFN__io_a_isInf = divSqrtRawFN_io_a_isSpecial & ~divSqrtRawFN_io_a_exp[21]; // @[rawFloatFromRecFN.scala 57:33]
  assign divSqrtRawFN__io_a_isZero = divSqrtRawFN_io_a_exp[23:21] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign divSqrtRawFN__io_a_sign = io_a[512]; // @[rawFloatFromRecFN.scala 59:25]
  assign divSqrtRawFN__io_a_sExp = {1'b0,$signed(divSqrtRawFN_io_a_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign divSqrtRawFN__io_a_sig = {_divSqrtRawFN_io_a_out_sig_T_1,io_a[487:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign divSqrtRawFN__io_b_isNaN = divSqrtRawFN_io_b_isSpecial & divSqrtRawFN_io_b_exp[21]; // @[rawFloatFromRecFN.scala 56:33]
  assign divSqrtRawFN__io_b_isInf = divSqrtRawFN_io_b_isSpecial & ~divSqrtRawFN_io_b_exp[21]; // @[rawFloatFromRecFN.scala 57:33]
  assign divSqrtRawFN__io_b_isZero = divSqrtRawFN_io_b_exp[23:21] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  assign divSqrtRawFN__io_b_sign = io_b[512]; // @[rawFloatFromRecFN.scala 59:25]
  assign divSqrtRawFN__io_b_sExp = {1'b0,$signed(divSqrtRawFN_io_b_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  assign divSqrtRawFN__io_b_sig = {_divSqrtRawFN_io_b_out_sig_T_1,io_b[487:0]}; // @[rawFloatFromRecFN.scala 61:44]
  assign divSqrtRawFN__io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 453:34]
endmodule
module RoundAnyRawFNToRecFN_ie23_is491_oe23_os489(
  input          io_invalidExc,
  input          io_infiniteExc,
  input          io_in_isNaN,
  input          io_in_isInf,
  input          io_in_isZero,
  input          io_in_sign,
  input  [24:0]  io_in_sExp,
  input  [491:0] io_in_sig,
  input  [2:0]   io_roundingMode,
  output [512:0] io_out,
  output [4:0]   io_exceptionFlags
);
  wire  roundingMode_near_even = io_roundingMode == 3'h0; // @[RoundAnyRawFNToRecFN.scala 90:53]
  wire  roundingMode_min = io_roundingMode == 3'h2; // @[RoundAnyRawFNToRecFN.scala 92:53]
  wire  roundingMode_max = io_roundingMode == 3'h3; // @[RoundAnyRawFNToRecFN.scala 93:53]
  wire  roundingMode_near_maxMag = io_roundingMode == 3'h4; // @[RoundAnyRawFNToRecFN.scala 94:53]
  wire  roundingMode_odd = io_roundingMode == 3'h6; // @[RoundAnyRawFNToRecFN.scala 95:53]
  wire  roundMagUp = roundingMode_min & io_in_sign | roundingMode_max & ~io_in_sign; // @[RoundAnyRawFNToRecFN.scala 98:42]
  wire  doShiftSigDown1 = io_in_sig[491]; // @[RoundAnyRawFNToRecFN.scala 120:57]
  wire [23:0] _roundMask_T_1 = ~io_in_sExp[23:0]; // @[primitives.scala 52:21]
  wire  roundMask_msb = _roundMask_T_1[23]; // @[primitives.scala 58:25]
  wire [22:0] roundMask_lsbs = _roundMask_T_1[22:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_1 = roundMask_lsbs[22]; // @[primitives.scala 58:25]
  wire [21:0] roundMask_lsbs_1 = roundMask_lsbs[21:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_2 = roundMask_lsbs_1[21]; // @[primitives.scala 58:25]
  wire [20:0] roundMask_lsbs_2 = roundMask_lsbs_1[20:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_3 = roundMask_lsbs_2[20]; // @[primitives.scala 58:25]
  wire [19:0] roundMask_lsbs_3 = roundMask_lsbs_2[19:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_4 = roundMask_lsbs_3[19]; // @[primitives.scala 58:25]
  wire [18:0] roundMask_lsbs_4 = roundMask_lsbs_3[18:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_5 = roundMask_lsbs_4[18]; // @[primitives.scala 58:25]
  wire [17:0] roundMask_lsbs_5 = roundMask_lsbs_4[17:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_6 = roundMask_lsbs_5[17]; // @[primitives.scala 58:25]
  wire [16:0] roundMask_lsbs_6 = roundMask_lsbs_5[16:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_7 = roundMask_lsbs_6[16]; // @[primitives.scala 58:25]
  wire [15:0] roundMask_lsbs_7 = roundMask_lsbs_6[15:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_8 = roundMask_lsbs_7[15]; // @[primitives.scala 58:25]
  wire [14:0] roundMask_lsbs_8 = roundMask_lsbs_7[14:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_9 = roundMask_lsbs_8[14]; // @[primitives.scala 58:25]
  wire [13:0] roundMask_lsbs_9 = roundMask_lsbs_8[13:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_10 = roundMask_lsbs_9[13]; // @[primitives.scala 58:25]
  wire [12:0] roundMask_lsbs_10 = roundMask_lsbs_9[12:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_11 = roundMask_lsbs_10[12]; // @[primitives.scala 58:25]
  wire [11:0] roundMask_lsbs_11 = roundMask_lsbs_10[11:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_12 = roundMask_lsbs_11[11]; // @[primitives.scala 58:25]
  wire [10:0] roundMask_lsbs_12 = roundMask_lsbs_11[10:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_13 = roundMask_lsbs_12[10]; // @[primitives.scala 58:25]
  wire [9:0] roundMask_lsbs_13 = roundMask_lsbs_12[9:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_14 = roundMask_lsbs_13[9]; // @[primitives.scala 58:25]
  wire [8:0] roundMask_lsbs_14 = roundMask_lsbs_13[8:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_15 = roundMask_lsbs_14[8]; // @[primitives.scala 58:25]
  wire [7:0] roundMask_lsbs_15 = roundMask_lsbs_14[7:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_16 = roundMask_lsbs_15[7]; // @[primitives.scala 58:25]
  wire [6:0] roundMask_lsbs_16 = roundMask_lsbs_15[6:0]; // @[primitives.scala 59:26]
  wire  roundMask_msb_17 = roundMask_lsbs_16[6]; // @[primitives.scala 58:25]
  wire [5:0] roundMask_lsbs_17 = roundMask_lsbs_16[5:0]; // @[primitives.scala 59:26]
  wire [64:0] roundMask_shift = 65'sh10000000000000000 >>> roundMask_lsbs_17; // @[primitives.scala 76:56]
  wire [31:0] _GEN_0 = {{16'd0}, roundMask_shift[56:41]}; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_7 = _GEN_0 & 32'hffff; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_9 = {roundMask_shift[40:25], 16'h0}; // @[Bitwise.scala 108:70]
  wire [31:0] _roundMask_T_11 = _roundMask_T_9 & 32'hffff0000; // @[Bitwise.scala 108:80]
  wire [31:0] _roundMask_T_12 = _roundMask_T_7 | _roundMask_T_11; // @[Bitwise.scala 108:39]
  wire [31:0] _GEN_1 = {{8'd0}, _roundMask_T_12[31:8]}; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_17 = _GEN_1 & 32'hff00ff; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_19 = {_roundMask_T_12[23:0], 8'h0}; // @[Bitwise.scala 108:70]
  wire [31:0] _roundMask_T_21 = _roundMask_T_19 & 32'hff00ff00; // @[Bitwise.scala 108:80]
  wire [31:0] _roundMask_T_22 = _roundMask_T_17 | _roundMask_T_21; // @[Bitwise.scala 108:39]
  wire [31:0] _GEN_2 = {{4'd0}, _roundMask_T_22[31:4]}; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_27 = _GEN_2 & 32'hf0f0f0f; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_29 = {_roundMask_T_22[27:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [31:0] _roundMask_T_31 = _roundMask_T_29 & 32'hf0f0f0f0; // @[Bitwise.scala 108:80]
  wire [31:0] _roundMask_T_32 = _roundMask_T_27 | _roundMask_T_31; // @[Bitwise.scala 108:39]
  wire [31:0] _GEN_3 = {{2'd0}, _roundMask_T_32[31:2]}; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_37 = _GEN_3 & 32'h33333333; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_39 = {_roundMask_T_32[29:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [31:0] _roundMask_T_41 = _roundMask_T_39 & 32'hcccccccc; // @[Bitwise.scala 108:80]
  wire [31:0] _roundMask_T_42 = _roundMask_T_37 | _roundMask_T_41; // @[Bitwise.scala 108:39]
  wire [31:0] _GEN_4 = {{1'd0}, _roundMask_T_42[31:1]}; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_47 = _GEN_4 & 32'h55555555; // @[Bitwise.scala 108:31]
  wire [31:0] _roundMask_T_49 = {_roundMask_T_42[30:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [31:0] _roundMask_T_51 = _roundMask_T_49 & 32'haaaaaaaa; // @[Bitwise.scala 108:80]
  wire [31:0] _roundMask_T_52 = _roundMask_T_47 | _roundMask_T_51; // @[Bitwise.scala 108:39]
  wire [102:0] _roundMask_T_73 = {_roundMask_T_52,roundMask_shift[57],roundMask_shift[58],roundMask_shift[59],
    roundMask_shift[60],roundMask_shift[61],roundMask_shift[62],roundMask_shift[63],64'hffffffffffffffff}; // @[primitives.scala 68:58]
  wire [63:0] _GEN_5 = {{32'd0}, roundMask_shift[63:32]}; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_78 = _GEN_5 & 64'hffffffff; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_80 = {roundMask_shift[31:0], 32'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _roundMask_T_82 = _roundMask_T_80 & 64'hffffffff00000000; // @[Bitwise.scala 108:80]
  wire [63:0] _roundMask_T_83 = _roundMask_T_78 | _roundMask_T_82; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_6 = {{16'd0}, _roundMask_T_83[63:16]}; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_88 = _GEN_6 & 64'hffff0000ffff; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_90 = {_roundMask_T_83[47:0], 16'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _roundMask_T_92 = _roundMask_T_90 & 64'hffff0000ffff0000; // @[Bitwise.scala 108:80]
  wire [63:0] _roundMask_T_93 = _roundMask_T_88 | _roundMask_T_92; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_7 = {{8'd0}, _roundMask_T_93[63:8]}; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_98 = _GEN_7 & 64'hff00ff00ff00ff; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_100 = {_roundMask_T_93[55:0], 8'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _roundMask_T_102 = _roundMask_T_100 & 64'hff00ff00ff00ff00; // @[Bitwise.scala 108:80]
  wire [63:0] _roundMask_T_103 = _roundMask_T_98 | _roundMask_T_102; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_8 = {{4'd0}, _roundMask_T_103[63:4]}; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_108 = _GEN_8 & 64'hf0f0f0f0f0f0f0f; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_110 = {_roundMask_T_103[59:0], 4'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _roundMask_T_112 = _roundMask_T_110 & 64'hf0f0f0f0f0f0f0f0; // @[Bitwise.scala 108:80]
  wire [63:0] _roundMask_T_113 = _roundMask_T_108 | _roundMask_T_112; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_9 = {{2'd0}, _roundMask_T_113[63:2]}; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_118 = _GEN_9 & 64'h3333333333333333; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_120 = {_roundMask_T_113[61:0], 2'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _roundMask_T_122 = _roundMask_T_120 & 64'hcccccccccccccccc; // @[Bitwise.scala 108:80]
  wire [63:0] _roundMask_T_123 = _roundMask_T_118 | _roundMask_T_122; // @[Bitwise.scala 108:39]
  wire [63:0] _GEN_10 = {{1'd0}, _roundMask_T_123[63:1]}; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_128 = _GEN_10 & 64'h5555555555555555; // @[Bitwise.scala 108:31]
  wire [63:0] _roundMask_T_130 = {_roundMask_T_123[62:0], 1'h0}; // @[Bitwise.scala 108:70]
  wire [63:0] _roundMask_T_132 = _roundMask_T_130 & 64'haaaaaaaaaaaaaaaa; // @[Bitwise.scala 108:80]
  wire [63:0] _roundMask_T_133 = _roundMask_T_128 | _roundMask_T_132; // @[Bitwise.scala 108:39]
  wire [102:0] _roundMask_T_134 = roundMask_msb_17 ? _roundMask_T_73 : {{39'd0}, _roundMask_T_133}; // @[primitives.scala 67:24]
  wire [230:0] _roundMask_T_135 = {_roundMask_T_134,128'hffffffffffffffffffffffffffffffff}; // @[primitives.scala 68:58]
  wire [127:0] _roundMask_T_196 = {_roundMask_T_133,64'hffffffffffffffff}; // @[primitives.scala 68:58]
  wire [127:0] _roundMask_T_257 = roundMask_msb_17 ? _roundMask_T_196 : {{64'd0}, _roundMask_T_133}; // @[primitives.scala 67:24]
  wire [230:0] _roundMask_T_258 = roundMask_msb_16 ? _roundMask_T_135 : {{103'd0}, _roundMask_T_257}; // @[primitives.scala 67:24]
  wire [486:0] _roundMask_T_259 = {_roundMask_T_258,256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
    }; // @[primitives.scala 68:58]
  wire [255:0] _roundMask_T_382 = {_roundMask_T_257,128'hffffffffffffffffffffffffffffffff}; // @[primitives.scala 68:58]
  wire [255:0] _roundMask_T_505 = roundMask_msb_16 ? _roundMask_T_382 : {{128'd0}, _roundMask_T_257}; // @[primitives.scala 67:24]
  wire [486:0] _roundMask_T_506 = roundMask_msb_15 ? _roundMask_T_259 : {{231'd0}, _roundMask_T_505}; // @[primitives.scala 67:24]
  wire [486:0] _roundMask_T_507 = ~_roundMask_T_506; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_508 = roundMask_msb_14 ? 487'h0 : _roundMask_T_507; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_509 = ~_roundMask_T_508; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_510 = ~_roundMask_T_509; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_511 = roundMask_msb_13 ? 487'h0 : _roundMask_T_510; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_512 = ~_roundMask_T_511; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_513 = ~_roundMask_T_512; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_514 = roundMask_msb_12 ? 487'h0 : _roundMask_T_513; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_515 = ~_roundMask_T_514; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_516 = ~_roundMask_T_515; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_517 = roundMask_msb_11 ? 487'h0 : _roundMask_T_516; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_518 = ~_roundMask_T_517; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_519 = ~_roundMask_T_518; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_520 = roundMask_msb_10 ? 487'h0 : _roundMask_T_519; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_521 = ~_roundMask_T_520; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_522 = ~_roundMask_T_521; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_523 = roundMask_msb_9 ? 487'h0 : _roundMask_T_522; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_524 = ~_roundMask_T_523; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_525 = ~_roundMask_T_524; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_526 = roundMask_msb_8 ? 487'h0 : _roundMask_T_525; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_527 = ~_roundMask_T_526; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_528 = ~_roundMask_T_527; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_529 = roundMask_msb_7 ? 487'h0 : _roundMask_T_528; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_530 = ~_roundMask_T_529; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_531 = ~_roundMask_T_530; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_532 = roundMask_msb_6 ? 487'h0 : _roundMask_T_531; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_533 = ~_roundMask_T_532; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_534 = ~_roundMask_T_533; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_535 = roundMask_msb_5 ? 487'h0 : _roundMask_T_534; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_536 = ~_roundMask_T_535; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_537 = ~_roundMask_T_536; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_538 = roundMask_msb_4 ? 487'h0 : _roundMask_T_537; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_539 = ~_roundMask_T_538; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_540 = ~_roundMask_T_539; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_541 = roundMask_msb_3 ? 487'h0 : _roundMask_T_540; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_542 = ~_roundMask_T_541; // @[primitives.scala 73:17]
  wire [486:0] _roundMask_T_543 = ~_roundMask_T_542; // @[primitives.scala 73:32]
  wire [486:0] _roundMask_T_544 = roundMask_msb_2 ? 487'h0 : _roundMask_T_543; // @[primitives.scala 73:21]
  wire [486:0] _roundMask_T_545 = ~_roundMask_T_544; // @[primitives.scala 73:17]
  wire [489:0] _roundMask_T_546 = {_roundMask_T_545,3'h7}; // @[primitives.scala 68:58]
  wire [2:0] _roundMask_T_553 = {roundMask_shift[0],roundMask_shift[1],roundMask_shift[2]}; // @[Cat.scala 33:92]
  wire [2:0] _roundMask_T_554 = roundMask_msb_17 ? _roundMask_T_553 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_555 = roundMask_msb_16 ? _roundMask_T_554 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_556 = roundMask_msb_15 ? _roundMask_T_555 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_557 = roundMask_msb_14 ? _roundMask_T_556 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_558 = roundMask_msb_13 ? _roundMask_T_557 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_559 = roundMask_msb_12 ? _roundMask_T_558 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_560 = roundMask_msb_11 ? _roundMask_T_559 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_561 = roundMask_msb_10 ? _roundMask_T_560 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_562 = roundMask_msb_9 ? _roundMask_T_561 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_563 = roundMask_msb_8 ? _roundMask_T_562 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_564 = roundMask_msb_7 ? _roundMask_T_563 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_565 = roundMask_msb_6 ? _roundMask_T_564 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_566 = roundMask_msb_5 ? _roundMask_T_565 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_567 = roundMask_msb_4 ? _roundMask_T_566 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_568 = roundMask_msb_3 ? _roundMask_T_567 : 3'h0; // @[primitives.scala 62:24]
  wire [2:0] _roundMask_T_569 = roundMask_msb_2 ? _roundMask_T_568 : 3'h0; // @[primitives.scala 62:24]
  wire [489:0] _roundMask_T_570 = roundMask_msb_1 ? _roundMask_T_546 : {{487'd0}, _roundMask_T_569}; // @[primitives.scala 67:24]
  wire [489:0] _roundMask_T_571 = roundMask_msb ? _roundMask_T_570 : 490'h0; // @[primitives.scala 62:24]
  wire [489:0] _GEN_47 = {{489'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 159:23]
  wire [489:0] _roundMask_T_572 = _roundMask_T_571 | _GEN_47; // @[RoundAnyRawFNToRecFN.scala 159:23]
  wire [491:0] roundMask = {_roundMask_T_572,2'h3}; // @[RoundAnyRawFNToRecFN.scala 159:42]
  wire [492:0] _shiftedRoundMask_T = {1'h0,_roundMask_T_572,2'h3}; // @[RoundAnyRawFNToRecFN.scala 162:41]
  wire [491:0] shiftedRoundMask = _shiftedRoundMask_T[492:1]; // @[RoundAnyRawFNToRecFN.scala 162:53]
  wire [491:0] _roundPosMask_T = ~shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 163:28]
  wire [491:0] roundPosMask = _roundPosMask_T & roundMask; // @[RoundAnyRawFNToRecFN.scala 163:46]
  wire [491:0] _roundPosBit_T = io_in_sig & roundPosMask; // @[RoundAnyRawFNToRecFN.scala 164:40]
  wire  roundPosBit = |_roundPosBit_T; // @[RoundAnyRawFNToRecFN.scala 164:56]
  wire [491:0] _anyRoundExtra_T = io_in_sig & shiftedRoundMask; // @[RoundAnyRawFNToRecFN.scala 165:42]
  wire  anyRoundExtra = |_anyRoundExtra_T; // @[RoundAnyRawFNToRecFN.scala 165:62]
  wire  anyRound = roundPosBit | anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 166:36]
  wire  _roundIncr_T = roundingMode_near_even | roundingMode_near_maxMag; // @[RoundAnyRawFNToRecFN.scala 169:38]
  wire  _roundIncr_T_1 = (roundingMode_near_even | roundingMode_near_maxMag) & roundPosBit; // @[RoundAnyRawFNToRecFN.scala 169:67]
  wire  _roundIncr_T_2 = roundMagUp & anyRound; // @[RoundAnyRawFNToRecFN.scala 171:29]
  wire  roundIncr = _roundIncr_T_1 | _roundIncr_T_2; // @[RoundAnyRawFNToRecFN.scala 170:31]
  wire [491:0] _roundedSig_T = io_in_sig | roundMask; // @[RoundAnyRawFNToRecFN.scala 174:32]
  wire [490:0] _roundedSig_T_2 = _roundedSig_T[491:2] + 490'h1; // @[RoundAnyRawFNToRecFN.scala 174:49]
  wire  _roundedSig_T_4 = ~anyRoundExtra; // @[RoundAnyRawFNToRecFN.scala 176:30]
  wire [490:0] _roundedSig_T_7 = roundingMode_near_even & roundPosBit & _roundedSig_T_4 ? roundMask[491:1] : 491'h0; // @[RoundAnyRawFNToRecFN.scala 175:25]
  wire [490:0] _roundedSig_T_8 = ~_roundedSig_T_7; // @[RoundAnyRawFNToRecFN.scala 175:21]
  wire [490:0] _roundedSig_T_9 = _roundedSig_T_2 & _roundedSig_T_8; // @[RoundAnyRawFNToRecFN.scala 174:57]
  wire [491:0] _roundedSig_T_10 = ~roundMask; // @[RoundAnyRawFNToRecFN.scala 180:32]
  wire [491:0] _roundedSig_T_11 = io_in_sig & _roundedSig_T_10; // @[RoundAnyRawFNToRecFN.scala 180:30]
  wire [490:0] _roundedSig_T_15 = roundingMode_odd & anyRound ? roundPosMask[491:1] : 491'h0; // @[RoundAnyRawFNToRecFN.scala 181:24]
  wire [490:0] _GEN_48 = {{1'd0}, _roundedSig_T_11[491:2]}; // @[RoundAnyRawFNToRecFN.scala 180:47]
  wire [490:0] _roundedSig_T_16 = _GEN_48 | _roundedSig_T_15; // @[RoundAnyRawFNToRecFN.scala 180:47]
  wire [490:0] roundedSig = roundIncr ? _roundedSig_T_9 : _roundedSig_T_16; // @[RoundAnyRawFNToRecFN.scala 173:16]
  wire [2:0] _sRoundedExp_T_1 = {1'b0,$signed(roundedSig[490:489])}; // @[RoundAnyRawFNToRecFN.scala 185:76]
  wire [24:0] _GEN_49 = {{22{_sRoundedExp_T_1[2]}},_sRoundedExp_T_1}; // @[RoundAnyRawFNToRecFN.scala 185:40]
  wire [25:0] sRoundedExp = $signed(io_in_sExp) + $signed(_GEN_49); // @[RoundAnyRawFNToRecFN.scala 185:40]
  wire [23:0] common_expOut = sRoundedExp[23:0]; // @[RoundAnyRawFNToRecFN.scala 187:37]
  wire [487:0] common_fractOut = doShiftSigDown1 ? roundedSig[488:1] : roundedSig[487:0]; // @[RoundAnyRawFNToRecFN.scala 189:16]
  wire [3:0] _common_overflow_T = sRoundedExp[25:22]; // @[RoundAnyRawFNToRecFN.scala 196:30]
  wire  common_overflow = $signed(_common_overflow_T) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 196:50]
  wire  common_totalUnderflow = $signed(sRoundedExp) < 26'sh3ffe1a; // @[RoundAnyRawFNToRecFN.scala 200:31]
  wire [1:0] _common_underflow_T = io_in_sExp[24:23]; // @[RoundAnyRawFNToRecFN.scala 220:49]
  wire  _common_underflow_T_5 = doShiftSigDown1 ? roundMask[3] : roundMask[2]; // @[RoundAnyRawFNToRecFN.scala 221:30]
  wire  _common_underflow_T_6 = anyRound & $signed(_common_underflow_T) <= 2'sh0 & _common_underflow_T_5; // @[RoundAnyRawFNToRecFN.scala 220:72]
  wire  common_underflow = common_totalUnderflow | _common_underflow_T_6; // @[RoundAnyRawFNToRecFN.scala 217:40]
  wire  common_inexact = common_totalUnderflow | anyRound; // @[RoundAnyRawFNToRecFN.scala 230:49]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 235:34]
  wire  notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 236:49]
  wire  commonCase = ~isNaNOut & ~notNaN_isSpecialInfOut & ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 237:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 238:32]
  wire  underflow = commonCase & common_underflow; // @[RoundAnyRawFNToRecFN.scala 239:32]
  wire  inexact = overflow | commonCase & common_inexact; // @[RoundAnyRawFNToRecFN.scala 240:28]
  wire  overflow_roundMagUp = _roundIncr_T | roundMagUp; // @[RoundAnyRawFNToRecFN.scala 243:60]
  wire  pegMinNonzeroMagOut = commonCase & common_totalUnderflow & (roundMagUp | roundingMode_odd); // @[RoundAnyRawFNToRecFN.scala 245:45]
  wire  pegMaxFiniteMagOut = overflow & ~overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 246:39]
  wire  notNaN_isInfOut = notNaN_isSpecialInfOut | overflow & overflow_roundMagUp; // @[RoundAnyRawFNToRecFN.scala 248:32]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 250:22]
  wire [23:0] _expOut_T_1 = io_in_isZero | common_totalUnderflow ? 24'he00000 : 24'h0; // @[RoundAnyRawFNToRecFN.scala 253:18]
  wire [23:0] _expOut_T_2 = ~_expOut_T_1; // @[RoundAnyRawFNToRecFN.scala 253:14]
  wire [23:0] _expOut_T_3 = common_expOut & _expOut_T_2; // @[RoundAnyRawFNToRecFN.scala 252:24]
  wire [23:0] _expOut_T_5 = pegMinNonzeroMagOut ? 24'hc001e5 : 24'h0; // @[RoundAnyRawFNToRecFN.scala 257:18]
  wire [23:0] _expOut_T_6 = ~_expOut_T_5; // @[RoundAnyRawFNToRecFN.scala 257:14]
  wire [23:0] _expOut_T_7 = _expOut_T_3 & _expOut_T_6; // @[RoundAnyRawFNToRecFN.scala 256:17]
  wire [23:0] _expOut_T_8 = pegMaxFiniteMagOut ? 24'h400000 : 24'h0; // @[RoundAnyRawFNToRecFN.scala 261:18]
  wire [23:0] _expOut_T_9 = ~_expOut_T_8; // @[RoundAnyRawFNToRecFN.scala 261:14]
  wire [23:0] _expOut_T_10 = _expOut_T_7 & _expOut_T_9; // @[RoundAnyRawFNToRecFN.scala 260:17]
  wire [23:0] _expOut_T_11 = notNaN_isInfOut ? 24'h200000 : 24'h0; // @[RoundAnyRawFNToRecFN.scala 265:18]
  wire [23:0] _expOut_T_12 = ~_expOut_T_11; // @[RoundAnyRawFNToRecFN.scala 265:14]
  wire [23:0] _expOut_T_13 = _expOut_T_10 & _expOut_T_12; // @[RoundAnyRawFNToRecFN.scala 264:17]
  wire [23:0] _expOut_T_14 = pegMinNonzeroMagOut ? 24'h3ffe1a : 24'h0; // @[RoundAnyRawFNToRecFN.scala 269:16]
  wire [23:0] _expOut_T_15 = _expOut_T_13 | _expOut_T_14; // @[RoundAnyRawFNToRecFN.scala 268:18]
  wire [23:0] _expOut_T_16 = pegMaxFiniteMagOut ? 24'hbfffff : 24'h0; // @[RoundAnyRawFNToRecFN.scala 273:16]
  wire [23:0] _expOut_T_17 = _expOut_T_15 | _expOut_T_16; // @[RoundAnyRawFNToRecFN.scala 272:15]
  wire [23:0] _expOut_T_18 = notNaN_isInfOut ? 24'hc00000 : 24'h0; // @[RoundAnyRawFNToRecFN.scala 277:16]
  wire [23:0] _expOut_T_19 = _expOut_T_17 | _expOut_T_18; // @[RoundAnyRawFNToRecFN.scala 276:15]
  wire [23:0] _expOut_T_20 = isNaNOut ? 24'he00000 : 24'h0; // @[RoundAnyRawFNToRecFN.scala 278:16]
  wire [23:0] expOut = _expOut_T_19 | _expOut_T_20; // @[RoundAnyRawFNToRecFN.scala 277:73]
  wire [487:0] _fractOut_T_2 = isNaNOut ? 488'h80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
     : 488'h0; // @[RoundAnyRawFNToRecFN.scala 281:16]
  wire [487:0] _fractOut_T_3 = isNaNOut | io_in_isZero | common_totalUnderflow ? _fractOut_T_2 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 280:12]
  wire [487:0] _fractOut_T_5 = pegMaxFiniteMagOut ? 488'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
     : 488'h0; // @[Bitwise.scala 77:12]
  wire [487:0] fractOut = _fractOut_T_3 | _fractOut_T_5; // @[RoundAnyRawFNToRecFN.scala 283:11]
  wire [24:0] _io_out_T = {signOut,expOut}; // @[RoundAnyRawFNToRecFN.scala 286:23]
  wire [3:0] _io_exceptionFlags_T_2 = {io_invalidExc,io_infiniteExc,overflow,underflow}; // @[RoundAnyRawFNToRecFN.scala 288:53]
  assign io_out = {_io_out_T,fractOut}; // @[RoundAnyRawFNToRecFN.scala 286:33]
  assign io_exceptionFlags = {_io_exceptionFlags_T_2,inexact}; // @[RoundAnyRawFNToRecFN.scala 288:66]
endmodule
module RoundRawFNToRecFN_e23_s489(
  input          io_invalidExc,
  input          io_infiniteExc,
  input          io_in_isNaN,
  input          io_in_isInf,
  input          io_in_isZero,
  input          io_in_sign,
  input  [24:0]  io_in_sExp,
  input  [491:0] io_in_sig,
  input  [2:0]   io_roundingMode,
  output [512:0] io_out,
  output [4:0]   io_exceptionFlags
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [24:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [491:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [2:0] roundAnyRawFNToRecFN_io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [512:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 310:15]
  wire [4:0] roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 310:15]
  RoundAnyRawFNToRecFN_ie23_is491_oe23_os489 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 310:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundAnyRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundAnyRawFNToRecFN_io_roundingMode),
    .io_out(roundAnyRawFNToRecFN_io_out),
    .io_exceptionFlags(roundAnyRawFNToRecFN_io_exceptionFlags)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 318:23]
  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags; // @[RoundAnyRawFNToRecFN.scala 319:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 313:44]
  assign roundAnyRawFNToRecFN_io_infiniteExc = io_infiniteExc; // @[RoundAnyRawFNToRecFN.scala 314:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 315:44]
  assign roundAnyRawFNToRecFN_io_roundingMode = io_roundingMode; // @[RoundAnyRawFNToRecFN.scala 316:44]
endmodule
module DivSqrtRecFM_small_e23_s489(
  input          clock,
  input          reset,
  output         io_inReady,
  input          io_inValid,
  input  [512:0] io_a,
  input  [512:0] io_b,
  input  [2:0]   io_roundingMode,
  output         io_outValid_div,
  output [512:0] io_out,
  output [4:0]   io_exceptionFlags
);
  wire  divSqrtRecFNToRaw_clock; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_reset; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_inValid; // @[DivSqrtRecFN_small.scala 493:15]
  wire [512:0] divSqrtRecFNToRaw_io_a; // @[DivSqrtRecFN_small.scala 493:15]
  wire [512:0] divSqrtRecFNToRaw_io_b; // @[DivSqrtRecFN_small.scala 493:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingMode; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 493:15]
  wire [2:0] divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 493:15]
  wire  divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 493:15]
  wire [24:0] divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 493:15]
  wire [491:0] divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 493:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[DivSqrtRecFN_small.scala 508:15]
  wire  roundRawFNToRecFN_io_infiniteExc; // @[DivSqrtRecFN_small.scala 508:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[DivSqrtRecFN_small.scala 508:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[DivSqrtRecFN_small.scala 508:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[DivSqrtRecFN_small.scala 508:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[DivSqrtRecFN_small.scala 508:15]
  wire [24:0] roundRawFNToRecFN_io_in_sExp; // @[DivSqrtRecFN_small.scala 508:15]
  wire [491:0] roundRawFNToRecFN_io_in_sig; // @[DivSqrtRecFN_small.scala 508:15]
  wire [2:0] roundRawFNToRecFN_io_roundingMode; // @[DivSqrtRecFN_small.scala 508:15]
  wire [512:0] roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 508:15]
  wire [4:0] roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 508:15]
  DivSqrtRecFMToRaw_small_e23_s489 divSqrtRecFNToRaw ( // @[DivSqrtRecFN_small.scala 493:15]
    .clock(divSqrtRecFNToRaw_clock),
    .reset(divSqrtRecFNToRaw_reset),
    .io_inReady(divSqrtRecFNToRaw_io_inReady),
    .io_inValid(divSqrtRecFNToRaw_io_inValid),
    .io_a(divSqrtRecFNToRaw_io_a),
    .io_b(divSqrtRecFNToRaw_io_b),
    .io_roundingMode(divSqrtRecFNToRaw_io_roundingMode),
    .io_rawOutValid_div(divSqrtRecFNToRaw_io_rawOutValid_div),
    .io_roundingModeOut(divSqrtRecFNToRaw_io_roundingModeOut),
    .io_invalidExc(divSqrtRecFNToRaw_io_invalidExc),
    .io_infiniteExc(divSqrtRecFNToRaw_io_infiniteExc),
    .io_rawOut_isNaN(divSqrtRecFNToRaw_io_rawOut_isNaN),
    .io_rawOut_isInf(divSqrtRecFNToRaw_io_rawOut_isInf),
    .io_rawOut_isZero(divSqrtRecFNToRaw_io_rawOut_isZero),
    .io_rawOut_sign(divSqrtRecFNToRaw_io_rawOut_sign),
    .io_rawOut_sExp(divSqrtRecFNToRaw_io_rawOut_sExp),
    .io_rawOut_sig(divSqrtRecFNToRaw_io_rawOut_sig)
  );
  RoundRawFNToRecFN_e23_s489 roundRawFNToRecFN ( // @[DivSqrtRecFN_small.scala 508:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_infiniteExc(roundRawFNToRecFN_io_infiniteExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_roundingMode(roundRawFNToRecFN_io_roundingMode),
    .io_out(roundRawFNToRecFN_io_out),
    .io_exceptionFlags(roundRawFNToRecFN_io_exceptionFlags)
  );
  assign io_inReady = divSqrtRecFNToRaw_io_inReady; // @[DivSqrtRecFN_small.scala 495:16]
  assign io_outValid_div = divSqrtRecFNToRaw_io_rawOutValid_div; // @[DivSqrtRecFN_small.scala 504:22]
  assign io_out = roundRawFNToRecFN_io_out; // @[DivSqrtRecFN_small.scala 514:23]
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags; // @[DivSqrtRecFN_small.scala 515:23]
  assign divSqrtRecFNToRaw_clock = clock;
  assign divSqrtRecFNToRaw_reset = reset;
  assign divSqrtRecFNToRaw_io_inValid = io_inValid; // @[DivSqrtRecFN_small.scala 496:39]
  assign divSqrtRecFNToRaw_io_a = io_a; // @[DivSqrtRecFN_small.scala 498:39]
  assign divSqrtRecFNToRaw_io_b = io_b; // @[DivSqrtRecFN_small.scala 499:39]
  assign divSqrtRecFNToRaw_io_roundingMode = io_roundingMode; // @[DivSqrtRecFN_small.scala 500:39]
  assign roundRawFNToRecFN_io_invalidExc = divSqrtRecFNToRaw_io_invalidExc; // @[DivSqrtRecFN_small.scala 509:39]
  assign roundRawFNToRecFN_io_infiniteExc = divSqrtRecFNToRaw_io_infiniteExc; // @[DivSqrtRecFN_small.scala 510:39]
  assign roundRawFNToRecFN_io_in_isNaN = divSqrtRecFNToRaw_io_rawOut_isNaN; // @[DivSqrtRecFN_small.scala 511:39]
  assign roundRawFNToRecFN_io_in_isInf = divSqrtRecFNToRaw_io_rawOut_isInf; // @[DivSqrtRecFN_small.scala 511:39]
  assign roundRawFNToRecFN_io_in_isZero = divSqrtRecFNToRaw_io_rawOut_isZero; // @[DivSqrtRecFN_small.scala 511:39]
  assign roundRawFNToRecFN_io_in_sign = divSqrtRecFNToRaw_io_rawOut_sign; // @[DivSqrtRecFN_small.scala 511:39]
  assign roundRawFNToRecFN_io_in_sExp = divSqrtRecFNToRaw_io_rawOut_sExp; // @[DivSqrtRecFN_small.scala 511:39]
  assign roundRawFNToRecFN_io_in_sig = divSqrtRecFNToRaw_io_rawOut_sig; // @[DivSqrtRecFN_small.scala 511:39]
  assign roundRawFNToRecFN_io_roundingMode = divSqrtRecFNToRaw_io_roundingModeOut; // @[DivSqrtRecFN_small.scala 512:39]
endmodule
module scientist(
  input          clock,
  input          reset,
  input          io_opSel,
  input  [511:0] io_a,
  input  [511:0] io_b,
  input  [511:0] io_c,
  input  [2:0]   io_roundingMode,
  output [511:0] io_out,
  output [4:0]   io_exceptionFlags
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  divsqrt_f0_clock; // @[Emitscientist.scala 39:26]
  wire  divsqrt_f0_reset; // @[Emitscientist.scala 39:26]
  wire  divsqrt_f0_io_inReady; // @[Emitscientist.scala 39:26]
  wire  divsqrt_f0_io_inValid; // @[Emitscientist.scala 39:26]
  wire [512:0] divsqrt_f0_io_a; // @[Emitscientist.scala 39:26]
  wire [512:0] divsqrt_f0_io_b; // @[Emitscientist.scala 39:26]
  wire [2:0] divsqrt_f0_io_roundingMode; // @[Emitscientist.scala 39:26]
  wire  divsqrt_f0_io_outValid_div; // @[Emitscientist.scala 39:26]
  wire [512:0] divsqrt_f0_io_out; // @[Emitscientist.scala 39:26]
  wire [4:0] divsqrt_f0_io_exceptionFlags; // @[Emitscientist.scala 39:26]
  wire  roundingMatches_0 = 3'h0 == io_roundingMode; // @[Emitscientist.scala 19:47]
  wire  fmt0_recA_rawIn_sign = io_a[511]; // @[rawFloatFromFN.scala 44:18]
  wire [22:0] fmt0_recA_rawIn_expIn = io_a[510:488]; // @[rawFloatFromFN.scala 45:19]
  wire [487:0] fmt0_recA_rawIn_fractIn = io_a[487:0]; // @[rawFloatFromFN.scala 46:21]
  wire  fmt0_recA_rawIn_isZeroExpIn = fmt0_recA_rawIn_expIn == 23'h0; // @[rawFloatFromFN.scala 48:30]
  wire  fmt0_recA_rawIn_isZeroFractIn = fmt0_recA_rawIn_fractIn == 488'h0; // @[rawFloatFromFN.scala 49:34]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_488 = fmt0_recA_rawIn_fractIn[1] ? 9'h1e6 : 9'h1e7; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_489 = fmt0_recA_rawIn_fractIn[2] ? 9'h1e5 : _fmt0_recA_rawIn_normDist_T_488; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_490 = fmt0_recA_rawIn_fractIn[3] ? 9'h1e4 : _fmt0_recA_rawIn_normDist_T_489; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_491 = fmt0_recA_rawIn_fractIn[4] ? 9'h1e3 : _fmt0_recA_rawIn_normDist_T_490; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_492 = fmt0_recA_rawIn_fractIn[5] ? 9'h1e2 : _fmt0_recA_rawIn_normDist_T_491; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_493 = fmt0_recA_rawIn_fractIn[6] ? 9'h1e1 : _fmt0_recA_rawIn_normDist_T_492; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_494 = fmt0_recA_rawIn_fractIn[7] ? 9'h1e0 : _fmt0_recA_rawIn_normDist_T_493; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_495 = fmt0_recA_rawIn_fractIn[8] ? 9'h1df : _fmt0_recA_rawIn_normDist_T_494; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_496 = fmt0_recA_rawIn_fractIn[9] ? 9'h1de : _fmt0_recA_rawIn_normDist_T_495; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_497 = fmt0_recA_rawIn_fractIn[10] ? 9'h1dd : _fmt0_recA_rawIn_normDist_T_496; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_498 = fmt0_recA_rawIn_fractIn[11] ? 9'h1dc : _fmt0_recA_rawIn_normDist_T_497; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_499 = fmt0_recA_rawIn_fractIn[12] ? 9'h1db : _fmt0_recA_rawIn_normDist_T_498; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_500 = fmt0_recA_rawIn_fractIn[13] ? 9'h1da : _fmt0_recA_rawIn_normDist_T_499; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_501 = fmt0_recA_rawIn_fractIn[14] ? 9'h1d9 : _fmt0_recA_rawIn_normDist_T_500; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_502 = fmt0_recA_rawIn_fractIn[15] ? 9'h1d8 : _fmt0_recA_rawIn_normDist_T_501; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_503 = fmt0_recA_rawIn_fractIn[16] ? 9'h1d7 : _fmt0_recA_rawIn_normDist_T_502; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_504 = fmt0_recA_rawIn_fractIn[17] ? 9'h1d6 : _fmt0_recA_rawIn_normDist_T_503; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_505 = fmt0_recA_rawIn_fractIn[18] ? 9'h1d5 : _fmt0_recA_rawIn_normDist_T_504; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_506 = fmt0_recA_rawIn_fractIn[19] ? 9'h1d4 : _fmt0_recA_rawIn_normDist_T_505; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_507 = fmt0_recA_rawIn_fractIn[20] ? 9'h1d3 : _fmt0_recA_rawIn_normDist_T_506; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_508 = fmt0_recA_rawIn_fractIn[21] ? 9'h1d2 : _fmt0_recA_rawIn_normDist_T_507; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_509 = fmt0_recA_rawIn_fractIn[22] ? 9'h1d1 : _fmt0_recA_rawIn_normDist_T_508; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_510 = fmt0_recA_rawIn_fractIn[23] ? 9'h1d0 : _fmt0_recA_rawIn_normDist_T_509; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_511 = fmt0_recA_rawIn_fractIn[24] ? 9'h1cf : _fmt0_recA_rawIn_normDist_T_510; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_512 = fmt0_recA_rawIn_fractIn[25] ? 9'h1ce : _fmt0_recA_rawIn_normDist_T_511; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_513 = fmt0_recA_rawIn_fractIn[26] ? 9'h1cd : _fmt0_recA_rawIn_normDist_T_512; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_514 = fmt0_recA_rawIn_fractIn[27] ? 9'h1cc : _fmt0_recA_rawIn_normDist_T_513; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_515 = fmt0_recA_rawIn_fractIn[28] ? 9'h1cb : _fmt0_recA_rawIn_normDist_T_514; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_516 = fmt0_recA_rawIn_fractIn[29] ? 9'h1ca : _fmt0_recA_rawIn_normDist_T_515; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_517 = fmt0_recA_rawIn_fractIn[30] ? 9'h1c9 : _fmt0_recA_rawIn_normDist_T_516; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_518 = fmt0_recA_rawIn_fractIn[31] ? 9'h1c8 : _fmt0_recA_rawIn_normDist_T_517; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_519 = fmt0_recA_rawIn_fractIn[32] ? 9'h1c7 : _fmt0_recA_rawIn_normDist_T_518; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_520 = fmt0_recA_rawIn_fractIn[33] ? 9'h1c6 : _fmt0_recA_rawIn_normDist_T_519; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_521 = fmt0_recA_rawIn_fractIn[34] ? 9'h1c5 : _fmt0_recA_rawIn_normDist_T_520; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_522 = fmt0_recA_rawIn_fractIn[35] ? 9'h1c4 : _fmt0_recA_rawIn_normDist_T_521; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_523 = fmt0_recA_rawIn_fractIn[36] ? 9'h1c3 : _fmt0_recA_rawIn_normDist_T_522; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_524 = fmt0_recA_rawIn_fractIn[37] ? 9'h1c2 : _fmt0_recA_rawIn_normDist_T_523; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_525 = fmt0_recA_rawIn_fractIn[38] ? 9'h1c1 : _fmt0_recA_rawIn_normDist_T_524; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_526 = fmt0_recA_rawIn_fractIn[39] ? 9'h1c0 : _fmt0_recA_rawIn_normDist_T_525; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_527 = fmt0_recA_rawIn_fractIn[40] ? 9'h1bf : _fmt0_recA_rawIn_normDist_T_526; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_528 = fmt0_recA_rawIn_fractIn[41] ? 9'h1be : _fmt0_recA_rawIn_normDist_T_527; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_529 = fmt0_recA_rawIn_fractIn[42] ? 9'h1bd : _fmt0_recA_rawIn_normDist_T_528; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_530 = fmt0_recA_rawIn_fractIn[43] ? 9'h1bc : _fmt0_recA_rawIn_normDist_T_529; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_531 = fmt0_recA_rawIn_fractIn[44] ? 9'h1bb : _fmt0_recA_rawIn_normDist_T_530; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_532 = fmt0_recA_rawIn_fractIn[45] ? 9'h1ba : _fmt0_recA_rawIn_normDist_T_531; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_533 = fmt0_recA_rawIn_fractIn[46] ? 9'h1b9 : _fmt0_recA_rawIn_normDist_T_532; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_534 = fmt0_recA_rawIn_fractIn[47] ? 9'h1b8 : _fmt0_recA_rawIn_normDist_T_533; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_535 = fmt0_recA_rawIn_fractIn[48] ? 9'h1b7 : _fmt0_recA_rawIn_normDist_T_534; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_536 = fmt0_recA_rawIn_fractIn[49] ? 9'h1b6 : _fmt0_recA_rawIn_normDist_T_535; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_537 = fmt0_recA_rawIn_fractIn[50] ? 9'h1b5 : _fmt0_recA_rawIn_normDist_T_536; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_538 = fmt0_recA_rawIn_fractIn[51] ? 9'h1b4 : _fmt0_recA_rawIn_normDist_T_537; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_539 = fmt0_recA_rawIn_fractIn[52] ? 9'h1b3 : _fmt0_recA_rawIn_normDist_T_538; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_540 = fmt0_recA_rawIn_fractIn[53] ? 9'h1b2 : _fmt0_recA_rawIn_normDist_T_539; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_541 = fmt0_recA_rawIn_fractIn[54] ? 9'h1b1 : _fmt0_recA_rawIn_normDist_T_540; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_542 = fmt0_recA_rawIn_fractIn[55] ? 9'h1b0 : _fmt0_recA_rawIn_normDist_T_541; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_543 = fmt0_recA_rawIn_fractIn[56] ? 9'h1af : _fmt0_recA_rawIn_normDist_T_542; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_544 = fmt0_recA_rawIn_fractIn[57] ? 9'h1ae : _fmt0_recA_rawIn_normDist_T_543; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_545 = fmt0_recA_rawIn_fractIn[58] ? 9'h1ad : _fmt0_recA_rawIn_normDist_T_544; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_546 = fmt0_recA_rawIn_fractIn[59] ? 9'h1ac : _fmt0_recA_rawIn_normDist_T_545; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_547 = fmt0_recA_rawIn_fractIn[60] ? 9'h1ab : _fmt0_recA_rawIn_normDist_T_546; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_548 = fmt0_recA_rawIn_fractIn[61] ? 9'h1aa : _fmt0_recA_rawIn_normDist_T_547; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_549 = fmt0_recA_rawIn_fractIn[62] ? 9'h1a9 : _fmt0_recA_rawIn_normDist_T_548; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_550 = fmt0_recA_rawIn_fractIn[63] ? 9'h1a8 : _fmt0_recA_rawIn_normDist_T_549; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_551 = fmt0_recA_rawIn_fractIn[64] ? 9'h1a7 : _fmt0_recA_rawIn_normDist_T_550; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_552 = fmt0_recA_rawIn_fractIn[65] ? 9'h1a6 : _fmt0_recA_rawIn_normDist_T_551; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_553 = fmt0_recA_rawIn_fractIn[66] ? 9'h1a5 : _fmt0_recA_rawIn_normDist_T_552; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_554 = fmt0_recA_rawIn_fractIn[67] ? 9'h1a4 : _fmt0_recA_rawIn_normDist_T_553; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_555 = fmt0_recA_rawIn_fractIn[68] ? 9'h1a3 : _fmt0_recA_rawIn_normDist_T_554; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_556 = fmt0_recA_rawIn_fractIn[69] ? 9'h1a2 : _fmt0_recA_rawIn_normDist_T_555; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_557 = fmt0_recA_rawIn_fractIn[70] ? 9'h1a1 : _fmt0_recA_rawIn_normDist_T_556; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_558 = fmt0_recA_rawIn_fractIn[71] ? 9'h1a0 : _fmt0_recA_rawIn_normDist_T_557; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_559 = fmt0_recA_rawIn_fractIn[72] ? 9'h19f : _fmt0_recA_rawIn_normDist_T_558; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_560 = fmt0_recA_rawIn_fractIn[73] ? 9'h19e : _fmt0_recA_rawIn_normDist_T_559; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_561 = fmt0_recA_rawIn_fractIn[74] ? 9'h19d : _fmt0_recA_rawIn_normDist_T_560; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_562 = fmt0_recA_rawIn_fractIn[75] ? 9'h19c : _fmt0_recA_rawIn_normDist_T_561; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_563 = fmt0_recA_rawIn_fractIn[76] ? 9'h19b : _fmt0_recA_rawIn_normDist_T_562; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_564 = fmt0_recA_rawIn_fractIn[77] ? 9'h19a : _fmt0_recA_rawIn_normDist_T_563; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_565 = fmt0_recA_rawIn_fractIn[78] ? 9'h199 : _fmt0_recA_rawIn_normDist_T_564; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_566 = fmt0_recA_rawIn_fractIn[79] ? 9'h198 : _fmt0_recA_rawIn_normDist_T_565; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_567 = fmt0_recA_rawIn_fractIn[80] ? 9'h197 : _fmt0_recA_rawIn_normDist_T_566; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_568 = fmt0_recA_rawIn_fractIn[81] ? 9'h196 : _fmt0_recA_rawIn_normDist_T_567; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_569 = fmt0_recA_rawIn_fractIn[82] ? 9'h195 : _fmt0_recA_rawIn_normDist_T_568; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_570 = fmt0_recA_rawIn_fractIn[83] ? 9'h194 : _fmt0_recA_rawIn_normDist_T_569; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_571 = fmt0_recA_rawIn_fractIn[84] ? 9'h193 : _fmt0_recA_rawIn_normDist_T_570; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_572 = fmt0_recA_rawIn_fractIn[85] ? 9'h192 : _fmt0_recA_rawIn_normDist_T_571; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_573 = fmt0_recA_rawIn_fractIn[86] ? 9'h191 : _fmt0_recA_rawIn_normDist_T_572; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_574 = fmt0_recA_rawIn_fractIn[87] ? 9'h190 : _fmt0_recA_rawIn_normDist_T_573; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_575 = fmt0_recA_rawIn_fractIn[88] ? 9'h18f : _fmt0_recA_rawIn_normDist_T_574; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_576 = fmt0_recA_rawIn_fractIn[89] ? 9'h18e : _fmt0_recA_rawIn_normDist_T_575; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_577 = fmt0_recA_rawIn_fractIn[90] ? 9'h18d : _fmt0_recA_rawIn_normDist_T_576; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_578 = fmt0_recA_rawIn_fractIn[91] ? 9'h18c : _fmt0_recA_rawIn_normDist_T_577; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_579 = fmt0_recA_rawIn_fractIn[92] ? 9'h18b : _fmt0_recA_rawIn_normDist_T_578; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_580 = fmt0_recA_rawIn_fractIn[93] ? 9'h18a : _fmt0_recA_rawIn_normDist_T_579; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_581 = fmt0_recA_rawIn_fractIn[94] ? 9'h189 : _fmt0_recA_rawIn_normDist_T_580; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_582 = fmt0_recA_rawIn_fractIn[95] ? 9'h188 : _fmt0_recA_rawIn_normDist_T_581; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_583 = fmt0_recA_rawIn_fractIn[96] ? 9'h187 : _fmt0_recA_rawIn_normDist_T_582; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_584 = fmt0_recA_rawIn_fractIn[97] ? 9'h186 : _fmt0_recA_rawIn_normDist_T_583; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_585 = fmt0_recA_rawIn_fractIn[98] ? 9'h185 : _fmt0_recA_rawIn_normDist_T_584; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_586 = fmt0_recA_rawIn_fractIn[99] ? 9'h184 : _fmt0_recA_rawIn_normDist_T_585; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_587 = fmt0_recA_rawIn_fractIn[100] ? 9'h183 : _fmt0_recA_rawIn_normDist_T_586; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_588 = fmt0_recA_rawIn_fractIn[101] ? 9'h182 : _fmt0_recA_rawIn_normDist_T_587; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_589 = fmt0_recA_rawIn_fractIn[102] ? 9'h181 : _fmt0_recA_rawIn_normDist_T_588; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_590 = fmt0_recA_rawIn_fractIn[103] ? 9'h180 : _fmt0_recA_rawIn_normDist_T_589; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_591 = fmt0_recA_rawIn_fractIn[104] ? 9'h17f : _fmt0_recA_rawIn_normDist_T_590; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_592 = fmt0_recA_rawIn_fractIn[105] ? 9'h17e : _fmt0_recA_rawIn_normDist_T_591; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_593 = fmt0_recA_rawIn_fractIn[106] ? 9'h17d : _fmt0_recA_rawIn_normDist_T_592; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_594 = fmt0_recA_rawIn_fractIn[107] ? 9'h17c : _fmt0_recA_rawIn_normDist_T_593; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_595 = fmt0_recA_rawIn_fractIn[108] ? 9'h17b : _fmt0_recA_rawIn_normDist_T_594; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_596 = fmt0_recA_rawIn_fractIn[109] ? 9'h17a : _fmt0_recA_rawIn_normDist_T_595; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_597 = fmt0_recA_rawIn_fractIn[110] ? 9'h179 : _fmt0_recA_rawIn_normDist_T_596; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_598 = fmt0_recA_rawIn_fractIn[111] ? 9'h178 : _fmt0_recA_rawIn_normDist_T_597; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_599 = fmt0_recA_rawIn_fractIn[112] ? 9'h177 : _fmt0_recA_rawIn_normDist_T_598; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_600 = fmt0_recA_rawIn_fractIn[113] ? 9'h176 : _fmt0_recA_rawIn_normDist_T_599; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_601 = fmt0_recA_rawIn_fractIn[114] ? 9'h175 : _fmt0_recA_rawIn_normDist_T_600; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_602 = fmt0_recA_rawIn_fractIn[115] ? 9'h174 : _fmt0_recA_rawIn_normDist_T_601; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_603 = fmt0_recA_rawIn_fractIn[116] ? 9'h173 : _fmt0_recA_rawIn_normDist_T_602; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_604 = fmt0_recA_rawIn_fractIn[117] ? 9'h172 : _fmt0_recA_rawIn_normDist_T_603; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_605 = fmt0_recA_rawIn_fractIn[118] ? 9'h171 : _fmt0_recA_rawIn_normDist_T_604; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_606 = fmt0_recA_rawIn_fractIn[119] ? 9'h170 : _fmt0_recA_rawIn_normDist_T_605; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_607 = fmt0_recA_rawIn_fractIn[120] ? 9'h16f : _fmt0_recA_rawIn_normDist_T_606; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_608 = fmt0_recA_rawIn_fractIn[121] ? 9'h16e : _fmt0_recA_rawIn_normDist_T_607; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_609 = fmt0_recA_rawIn_fractIn[122] ? 9'h16d : _fmt0_recA_rawIn_normDist_T_608; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_610 = fmt0_recA_rawIn_fractIn[123] ? 9'h16c : _fmt0_recA_rawIn_normDist_T_609; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_611 = fmt0_recA_rawIn_fractIn[124] ? 9'h16b : _fmt0_recA_rawIn_normDist_T_610; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_612 = fmt0_recA_rawIn_fractIn[125] ? 9'h16a : _fmt0_recA_rawIn_normDist_T_611; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_613 = fmt0_recA_rawIn_fractIn[126] ? 9'h169 : _fmt0_recA_rawIn_normDist_T_612; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_614 = fmt0_recA_rawIn_fractIn[127] ? 9'h168 : _fmt0_recA_rawIn_normDist_T_613; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_615 = fmt0_recA_rawIn_fractIn[128] ? 9'h167 : _fmt0_recA_rawIn_normDist_T_614; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_616 = fmt0_recA_rawIn_fractIn[129] ? 9'h166 : _fmt0_recA_rawIn_normDist_T_615; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_617 = fmt0_recA_rawIn_fractIn[130] ? 9'h165 : _fmt0_recA_rawIn_normDist_T_616; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_618 = fmt0_recA_rawIn_fractIn[131] ? 9'h164 : _fmt0_recA_rawIn_normDist_T_617; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_619 = fmt0_recA_rawIn_fractIn[132] ? 9'h163 : _fmt0_recA_rawIn_normDist_T_618; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_620 = fmt0_recA_rawIn_fractIn[133] ? 9'h162 : _fmt0_recA_rawIn_normDist_T_619; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_621 = fmt0_recA_rawIn_fractIn[134] ? 9'h161 : _fmt0_recA_rawIn_normDist_T_620; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_622 = fmt0_recA_rawIn_fractIn[135] ? 9'h160 : _fmt0_recA_rawIn_normDist_T_621; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_623 = fmt0_recA_rawIn_fractIn[136] ? 9'h15f : _fmt0_recA_rawIn_normDist_T_622; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_624 = fmt0_recA_rawIn_fractIn[137] ? 9'h15e : _fmt0_recA_rawIn_normDist_T_623; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_625 = fmt0_recA_rawIn_fractIn[138] ? 9'h15d : _fmt0_recA_rawIn_normDist_T_624; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_626 = fmt0_recA_rawIn_fractIn[139] ? 9'h15c : _fmt0_recA_rawIn_normDist_T_625; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_627 = fmt0_recA_rawIn_fractIn[140] ? 9'h15b : _fmt0_recA_rawIn_normDist_T_626; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_628 = fmt0_recA_rawIn_fractIn[141] ? 9'h15a : _fmt0_recA_rawIn_normDist_T_627; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_629 = fmt0_recA_rawIn_fractIn[142] ? 9'h159 : _fmt0_recA_rawIn_normDist_T_628; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_630 = fmt0_recA_rawIn_fractIn[143] ? 9'h158 : _fmt0_recA_rawIn_normDist_T_629; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_631 = fmt0_recA_rawIn_fractIn[144] ? 9'h157 : _fmt0_recA_rawIn_normDist_T_630; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_632 = fmt0_recA_rawIn_fractIn[145] ? 9'h156 : _fmt0_recA_rawIn_normDist_T_631; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_633 = fmt0_recA_rawIn_fractIn[146] ? 9'h155 : _fmt0_recA_rawIn_normDist_T_632; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_634 = fmt0_recA_rawIn_fractIn[147] ? 9'h154 : _fmt0_recA_rawIn_normDist_T_633; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_635 = fmt0_recA_rawIn_fractIn[148] ? 9'h153 : _fmt0_recA_rawIn_normDist_T_634; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_636 = fmt0_recA_rawIn_fractIn[149] ? 9'h152 : _fmt0_recA_rawIn_normDist_T_635; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_637 = fmt0_recA_rawIn_fractIn[150] ? 9'h151 : _fmt0_recA_rawIn_normDist_T_636; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_638 = fmt0_recA_rawIn_fractIn[151] ? 9'h150 : _fmt0_recA_rawIn_normDist_T_637; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_639 = fmt0_recA_rawIn_fractIn[152] ? 9'h14f : _fmt0_recA_rawIn_normDist_T_638; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_640 = fmt0_recA_rawIn_fractIn[153] ? 9'h14e : _fmt0_recA_rawIn_normDist_T_639; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_641 = fmt0_recA_rawIn_fractIn[154] ? 9'h14d : _fmt0_recA_rawIn_normDist_T_640; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_642 = fmt0_recA_rawIn_fractIn[155] ? 9'h14c : _fmt0_recA_rawIn_normDist_T_641; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_643 = fmt0_recA_rawIn_fractIn[156] ? 9'h14b : _fmt0_recA_rawIn_normDist_T_642; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_644 = fmt0_recA_rawIn_fractIn[157] ? 9'h14a : _fmt0_recA_rawIn_normDist_T_643; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_645 = fmt0_recA_rawIn_fractIn[158] ? 9'h149 : _fmt0_recA_rawIn_normDist_T_644; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_646 = fmt0_recA_rawIn_fractIn[159] ? 9'h148 : _fmt0_recA_rawIn_normDist_T_645; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_647 = fmt0_recA_rawIn_fractIn[160] ? 9'h147 : _fmt0_recA_rawIn_normDist_T_646; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_648 = fmt0_recA_rawIn_fractIn[161] ? 9'h146 : _fmt0_recA_rawIn_normDist_T_647; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_649 = fmt0_recA_rawIn_fractIn[162] ? 9'h145 : _fmt0_recA_rawIn_normDist_T_648; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_650 = fmt0_recA_rawIn_fractIn[163] ? 9'h144 : _fmt0_recA_rawIn_normDist_T_649; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_651 = fmt0_recA_rawIn_fractIn[164] ? 9'h143 : _fmt0_recA_rawIn_normDist_T_650; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_652 = fmt0_recA_rawIn_fractIn[165] ? 9'h142 : _fmt0_recA_rawIn_normDist_T_651; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_653 = fmt0_recA_rawIn_fractIn[166] ? 9'h141 : _fmt0_recA_rawIn_normDist_T_652; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_654 = fmt0_recA_rawIn_fractIn[167] ? 9'h140 : _fmt0_recA_rawIn_normDist_T_653; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_655 = fmt0_recA_rawIn_fractIn[168] ? 9'h13f : _fmt0_recA_rawIn_normDist_T_654; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_656 = fmt0_recA_rawIn_fractIn[169] ? 9'h13e : _fmt0_recA_rawIn_normDist_T_655; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_657 = fmt0_recA_rawIn_fractIn[170] ? 9'h13d : _fmt0_recA_rawIn_normDist_T_656; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_658 = fmt0_recA_rawIn_fractIn[171] ? 9'h13c : _fmt0_recA_rawIn_normDist_T_657; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_659 = fmt0_recA_rawIn_fractIn[172] ? 9'h13b : _fmt0_recA_rawIn_normDist_T_658; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_660 = fmt0_recA_rawIn_fractIn[173] ? 9'h13a : _fmt0_recA_rawIn_normDist_T_659; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_661 = fmt0_recA_rawIn_fractIn[174] ? 9'h139 : _fmt0_recA_rawIn_normDist_T_660; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_662 = fmt0_recA_rawIn_fractIn[175] ? 9'h138 : _fmt0_recA_rawIn_normDist_T_661; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_663 = fmt0_recA_rawIn_fractIn[176] ? 9'h137 : _fmt0_recA_rawIn_normDist_T_662; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_664 = fmt0_recA_rawIn_fractIn[177] ? 9'h136 : _fmt0_recA_rawIn_normDist_T_663; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_665 = fmt0_recA_rawIn_fractIn[178] ? 9'h135 : _fmt0_recA_rawIn_normDist_T_664; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_666 = fmt0_recA_rawIn_fractIn[179] ? 9'h134 : _fmt0_recA_rawIn_normDist_T_665; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_667 = fmt0_recA_rawIn_fractIn[180] ? 9'h133 : _fmt0_recA_rawIn_normDist_T_666; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_668 = fmt0_recA_rawIn_fractIn[181] ? 9'h132 : _fmt0_recA_rawIn_normDist_T_667; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_669 = fmt0_recA_rawIn_fractIn[182] ? 9'h131 : _fmt0_recA_rawIn_normDist_T_668; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_670 = fmt0_recA_rawIn_fractIn[183] ? 9'h130 : _fmt0_recA_rawIn_normDist_T_669; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_671 = fmt0_recA_rawIn_fractIn[184] ? 9'h12f : _fmt0_recA_rawIn_normDist_T_670; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_672 = fmt0_recA_rawIn_fractIn[185] ? 9'h12e : _fmt0_recA_rawIn_normDist_T_671; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_673 = fmt0_recA_rawIn_fractIn[186] ? 9'h12d : _fmt0_recA_rawIn_normDist_T_672; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_674 = fmt0_recA_rawIn_fractIn[187] ? 9'h12c : _fmt0_recA_rawIn_normDist_T_673; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_675 = fmt0_recA_rawIn_fractIn[188] ? 9'h12b : _fmt0_recA_rawIn_normDist_T_674; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_676 = fmt0_recA_rawIn_fractIn[189] ? 9'h12a : _fmt0_recA_rawIn_normDist_T_675; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_677 = fmt0_recA_rawIn_fractIn[190] ? 9'h129 : _fmt0_recA_rawIn_normDist_T_676; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_678 = fmt0_recA_rawIn_fractIn[191] ? 9'h128 : _fmt0_recA_rawIn_normDist_T_677; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_679 = fmt0_recA_rawIn_fractIn[192] ? 9'h127 : _fmt0_recA_rawIn_normDist_T_678; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_680 = fmt0_recA_rawIn_fractIn[193] ? 9'h126 : _fmt0_recA_rawIn_normDist_T_679; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_681 = fmt0_recA_rawIn_fractIn[194] ? 9'h125 : _fmt0_recA_rawIn_normDist_T_680; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_682 = fmt0_recA_rawIn_fractIn[195] ? 9'h124 : _fmt0_recA_rawIn_normDist_T_681; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_683 = fmt0_recA_rawIn_fractIn[196] ? 9'h123 : _fmt0_recA_rawIn_normDist_T_682; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_684 = fmt0_recA_rawIn_fractIn[197] ? 9'h122 : _fmt0_recA_rawIn_normDist_T_683; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_685 = fmt0_recA_rawIn_fractIn[198] ? 9'h121 : _fmt0_recA_rawIn_normDist_T_684; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_686 = fmt0_recA_rawIn_fractIn[199] ? 9'h120 : _fmt0_recA_rawIn_normDist_T_685; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_687 = fmt0_recA_rawIn_fractIn[200] ? 9'h11f : _fmt0_recA_rawIn_normDist_T_686; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_688 = fmt0_recA_rawIn_fractIn[201] ? 9'h11e : _fmt0_recA_rawIn_normDist_T_687; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_689 = fmt0_recA_rawIn_fractIn[202] ? 9'h11d : _fmt0_recA_rawIn_normDist_T_688; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_690 = fmt0_recA_rawIn_fractIn[203] ? 9'h11c : _fmt0_recA_rawIn_normDist_T_689; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_691 = fmt0_recA_rawIn_fractIn[204] ? 9'h11b : _fmt0_recA_rawIn_normDist_T_690; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_692 = fmt0_recA_rawIn_fractIn[205] ? 9'h11a : _fmt0_recA_rawIn_normDist_T_691; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_693 = fmt0_recA_rawIn_fractIn[206] ? 9'h119 : _fmt0_recA_rawIn_normDist_T_692; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_694 = fmt0_recA_rawIn_fractIn[207] ? 9'h118 : _fmt0_recA_rawIn_normDist_T_693; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_695 = fmt0_recA_rawIn_fractIn[208] ? 9'h117 : _fmt0_recA_rawIn_normDist_T_694; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_696 = fmt0_recA_rawIn_fractIn[209] ? 9'h116 : _fmt0_recA_rawIn_normDist_T_695; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_697 = fmt0_recA_rawIn_fractIn[210] ? 9'h115 : _fmt0_recA_rawIn_normDist_T_696; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_698 = fmt0_recA_rawIn_fractIn[211] ? 9'h114 : _fmt0_recA_rawIn_normDist_T_697; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_699 = fmt0_recA_rawIn_fractIn[212] ? 9'h113 : _fmt0_recA_rawIn_normDist_T_698; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_700 = fmt0_recA_rawIn_fractIn[213] ? 9'h112 : _fmt0_recA_rawIn_normDist_T_699; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_701 = fmt0_recA_rawIn_fractIn[214] ? 9'h111 : _fmt0_recA_rawIn_normDist_T_700; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_702 = fmt0_recA_rawIn_fractIn[215] ? 9'h110 : _fmt0_recA_rawIn_normDist_T_701; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_703 = fmt0_recA_rawIn_fractIn[216] ? 9'h10f : _fmt0_recA_rawIn_normDist_T_702; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_704 = fmt0_recA_rawIn_fractIn[217] ? 9'h10e : _fmt0_recA_rawIn_normDist_T_703; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_705 = fmt0_recA_rawIn_fractIn[218] ? 9'h10d : _fmt0_recA_rawIn_normDist_T_704; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_706 = fmt0_recA_rawIn_fractIn[219] ? 9'h10c : _fmt0_recA_rawIn_normDist_T_705; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_707 = fmt0_recA_rawIn_fractIn[220] ? 9'h10b : _fmt0_recA_rawIn_normDist_T_706; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_708 = fmt0_recA_rawIn_fractIn[221] ? 9'h10a : _fmt0_recA_rawIn_normDist_T_707; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_709 = fmt0_recA_rawIn_fractIn[222] ? 9'h109 : _fmt0_recA_rawIn_normDist_T_708; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_710 = fmt0_recA_rawIn_fractIn[223] ? 9'h108 : _fmt0_recA_rawIn_normDist_T_709; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_711 = fmt0_recA_rawIn_fractIn[224] ? 9'h107 : _fmt0_recA_rawIn_normDist_T_710; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_712 = fmt0_recA_rawIn_fractIn[225] ? 9'h106 : _fmt0_recA_rawIn_normDist_T_711; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_713 = fmt0_recA_rawIn_fractIn[226] ? 9'h105 : _fmt0_recA_rawIn_normDist_T_712; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_714 = fmt0_recA_rawIn_fractIn[227] ? 9'h104 : _fmt0_recA_rawIn_normDist_T_713; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_715 = fmt0_recA_rawIn_fractIn[228] ? 9'h103 : _fmt0_recA_rawIn_normDist_T_714; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_716 = fmt0_recA_rawIn_fractIn[229] ? 9'h102 : _fmt0_recA_rawIn_normDist_T_715; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_717 = fmt0_recA_rawIn_fractIn[230] ? 9'h101 : _fmt0_recA_rawIn_normDist_T_716; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_718 = fmt0_recA_rawIn_fractIn[231] ? 9'h100 : _fmt0_recA_rawIn_normDist_T_717; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_719 = fmt0_recA_rawIn_fractIn[232] ? 9'hff : _fmt0_recA_rawIn_normDist_T_718; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_720 = fmt0_recA_rawIn_fractIn[233] ? 9'hfe : _fmt0_recA_rawIn_normDist_T_719; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_721 = fmt0_recA_rawIn_fractIn[234] ? 9'hfd : _fmt0_recA_rawIn_normDist_T_720; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_722 = fmt0_recA_rawIn_fractIn[235] ? 9'hfc : _fmt0_recA_rawIn_normDist_T_721; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_723 = fmt0_recA_rawIn_fractIn[236] ? 9'hfb : _fmt0_recA_rawIn_normDist_T_722; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_724 = fmt0_recA_rawIn_fractIn[237] ? 9'hfa : _fmt0_recA_rawIn_normDist_T_723; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_725 = fmt0_recA_rawIn_fractIn[238] ? 9'hf9 : _fmt0_recA_rawIn_normDist_T_724; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_726 = fmt0_recA_rawIn_fractIn[239] ? 9'hf8 : _fmt0_recA_rawIn_normDist_T_725; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_727 = fmt0_recA_rawIn_fractIn[240] ? 9'hf7 : _fmt0_recA_rawIn_normDist_T_726; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_728 = fmt0_recA_rawIn_fractIn[241] ? 9'hf6 : _fmt0_recA_rawIn_normDist_T_727; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_729 = fmt0_recA_rawIn_fractIn[242] ? 9'hf5 : _fmt0_recA_rawIn_normDist_T_728; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_730 = fmt0_recA_rawIn_fractIn[243] ? 9'hf4 : _fmt0_recA_rawIn_normDist_T_729; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_731 = fmt0_recA_rawIn_fractIn[244] ? 9'hf3 : _fmt0_recA_rawIn_normDist_T_730; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_732 = fmt0_recA_rawIn_fractIn[245] ? 9'hf2 : _fmt0_recA_rawIn_normDist_T_731; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_733 = fmt0_recA_rawIn_fractIn[246] ? 9'hf1 : _fmt0_recA_rawIn_normDist_T_732; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_734 = fmt0_recA_rawIn_fractIn[247] ? 9'hf0 : _fmt0_recA_rawIn_normDist_T_733; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_735 = fmt0_recA_rawIn_fractIn[248] ? 9'hef : _fmt0_recA_rawIn_normDist_T_734; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_736 = fmt0_recA_rawIn_fractIn[249] ? 9'hee : _fmt0_recA_rawIn_normDist_T_735; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_737 = fmt0_recA_rawIn_fractIn[250] ? 9'hed : _fmt0_recA_rawIn_normDist_T_736; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_738 = fmt0_recA_rawIn_fractIn[251] ? 9'hec : _fmt0_recA_rawIn_normDist_T_737; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_739 = fmt0_recA_rawIn_fractIn[252] ? 9'heb : _fmt0_recA_rawIn_normDist_T_738; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_740 = fmt0_recA_rawIn_fractIn[253] ? 9'hea : _fmt0_recA_rawIn_normDist_T_739; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_741 = fmt0_recA_rawIn_fractIn[254] ? 9'he9 : _fmt0_recA_rawIn_normDist_T_740; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_742 = fmt0_recA_rawIn_fractIn[255] ? 9'he8 : _fmt0_recA_rawIn_normDist_T_741; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_743 = fmt0_recA_rawIn_fractIn[256] ? 9'he7 : _fmt0_recA_rawIn_normDist_T_742; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_744 = fmt0_recA_rawIn_fractIn[257] ? 9'he6 : _fmt0_recA_rawIn_normDist_T_743; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_745 = fmt0_recA_rawIn_fractIn[258] ? 9'he5 : _fmt0_recA_rawIn_normDist_T_744; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_746 = fmt0_recA_rawIn_fractIn[259] ? 9'he4 : _fmt0_recA_rawIn_normDist_T_745; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_747 = fmt0_recA_rawIn_fractIn[260] ? 9'he3 : _fmt0_recA_rawIn_normDist_T_746; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_748 = fmt0_recA_rawIn_fractIn[261] ? 9'he2 : _fmt0_recA_rawIn_normDist_T_747; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_749 = fmt0_recA_rawIn_fractIn[262] ? 9'he1 : _fmt0_recA_rawIn_normDist_T_748; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_750 = fmt0_recA_rawIn_fractIn[263] ? 9'he0 : _fmt0_recA_rawIn_normDist_T_749; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_751 = fmt0_recA_rawIn_fractIn[264] ? 9'hdf : _fmt0_recA_rawIn_normDist_T_750; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_752 = fmt0_recA_rawIn_fractIn[265] ? 9'hde : _fmt0_recA_rawIn_normDist_T_751; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_753 = fmt0_recA_rawIn_fractIn[266] ? 9'hdd : _fmt0_recA_rawIn_normDist_T_752; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_754 = fmt0_recA_rawIn_fractIn[267] ? 9'hdc : _fmt0_recA_rawIn_normDist_T_753; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_755 = fmt0_recA_rawIn_fractIn[268] ? 9'hdb : _fmt0_recA_rawIn_normDist_T_754; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_756 = fmt0_recA_rawIn_fractIn[269] ? 9'hda : _fmt0_recA_rawIn_normDist_T_755; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_757 = fmt0_recA_rawIn_fractIn[270] ? 9'hd9 : _fmt0_recA_rawIn_normDist_T_756; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_758 = fmt0_recA_rawIn_fractIn[271] ? 9'hd8 : _fmt0_recA_rawIn_normDist_T_757; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_759 = fmt0_recA_rawIn_fractIn[272] ? 9'hd7 : _fmt0_recA_rawIn_normDist_T_758; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_760 = fmt0_recA_rawIn_fractIn[273] ? 9'hd6 : _fmt0_recA_rawIn_normDist_T_759; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_761 = fmt0_recA_rawIn_fractIn[274] ? 9'hd5 : _fmt0_recA_rawIn_normDist_T_760; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_762 = fmt0_recA_rawIn_fractIn[275] ? 9'hd4 : _fmt0_recA_rawIn_normDist_T_761; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_763 = fmt0_recA_rawIn_fractIn[276] ? 9'hd3 : _fmt0_recA_rawIn_normDist_T_762; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_764 = fmt0_recA_rawIn_fractIn[277] ? 9'hd2 : _fmt0_recA_rawIn_normDist_T_763; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_765 = fmt0_recA_rawIn_fractIn[278] ? 9'hd1 : _fmt0_recA_rawIn_normDist_T_764; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_766 = fmt0_recA_rawIn_fractIn[279] ? 9'hd0 : _fmt0_recA_rawIn_normDist_T_765; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_767 = fmt0_recA_rawIn_fractIn[280] ? 9'hcf : _fmt0_recA_rawIn_normDist_T_766; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_768 = fmt0_recA_rawIn_fractIn[281] ? 9'hce : _fmt0_recA_rawIn_normDist_T_767; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_769 = fmt0_recA_rawIn_fractIn[282] ? 9'hcd : _fmt0_recA_rawIn_normDist_T_768; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_770 = fmt0_recA_rawIn_fractIn[283] ? 9'hcc : _fmt0_recA_rawIn_normDist_T_769; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_771 = fmt0_recA_rawIn_fractIn[284] ? 9'hcb : _fmt0_recA_rawIn_normDist_T_770; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_772 = fmt0_recA_rawIn_fractIn[285] ? 9'hca : _fmt0_recA_rawIn_normDist_T_771; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_773 = fmt0_recA_rawIn_fractIn[286] ? 9'hc9 : _fmt0_recA_rawIn_normDist_T_772; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_774 = fmt0_recA_rawIn_fractIn[287] ? 9'hc8 : _fmt0_recA_rawIn_normDist_T_773; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_775 = fmt0_recA_rawIn_fractIn[288] ? 9'hc7 : _fmt0_recA_rawIn_normDist_T_774; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_776 = fmt0_recA_rawIn_fractIn[289] ? 9'hc6 : _fmt0_recA_rawIn_normDist_T_775; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_777 = fmt0_recA_rawIn_fractIn[290] ? 9'hc5 : _fmt0_recA_rawIn_normDist_T_776; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_778 = fmt0_recA_rawIn_fractIn[291] ? 9'hc4 : _fmt0_recA_rawIn_normDist_T_777; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_779 = fmt0_recA_rawIn_fractIn[292] ? 9'hc3 : _fmt0_recA_rawIn_normDist_T_778; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_780 = fmt0_recA_rawIn_fractIn[293] ? 9'hc2 : _fmt0_recA_rawIn_normDist_T_779; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_781 = fmt0_recA_rawIn_fractIn[294] ? 9'hc1 : _fmt0_recA_rawIn_normDist_T_780; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_782 = fmt0_recA_rawIn_fractIn[295] ? 9'hc0 : _fmt0_recA_rawIn_normDist_T_781; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_783 = fmt0_recA_rawIn_fractIn[296] ? 9'hbf : _fmt0_recA_rawIn_normDist_T_782; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_784 = fmt0_recA_rawIn_fractIn[297] ? 9'hbe : _fmt0_recA_rawIn_normDist_T_783; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_785 = fmt0_recA_rawIn_fractIn[298] ? 9'hbd : _fmt0_recA_rawIn_normDist_T_784; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_786 = fmt0_recA_rawIn_fractIn[299] ? 9'hbc : _fmt0_recA_rawIn_normDist_T_785; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_787 = fmt0_recA_rawIn_fractIn[300] ? 9'hbb : _fmt0_recA_rawIn_normDist_T_786; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_788 = fmt0_recA_rawIn_fractIn[301] ? 9'hba : _fmt0_recA_rawIn_normDist_T_787; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_789 = fmt0_recA_rawIn_fractIn[302] ? 9'hb9 : _fmt0_recA_rawIn_normDist_T_788; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_790 = fmt0_recA_rawIn_fractIn[303] ? 9'hb8 : _fmt0_recA_rawIn_normDist_T_789; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_791 = fmt0_recA_rawIn_fractIn[304] ? 9'hb7 : _fmt0_recA_rawIn_normDist_T_790; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_792 = fmt0_recA_rawIn_fractIn[305] ? 9'hb6 : _fmt0_recA_rawIn_normDist_T_791; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_793 = fmt0_recA_rawIn_fractIn[306] ? 9'hb5 : _fmt0_recA_rawIn_normDist_T_792; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_794 = fmt0_recA_rawIn_fractIn[307] ? 9'hb4 : _fmt0_recA_rawIn_normDist_T_793; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_795 = fmt0_recA_rawIn_fractIn[308] ? 9'hb3 : _fmt0_recA_rawIn_normDist_T_794; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_796 = fmt0_recA_rawIn_fractIn[309] ? 9'hb2 : _fmt0_recA_rawIn_normDist_T_795; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_797 = fmt0_recA_rawIn_fractIn[310] ? 9'hb1 : _fmt0_recA_rawIn_normDist_T_796; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_798 = fmt0_recA_rawIn_fractIn[311] ? 9'hb0 : _fmt0_recA_rawIn_normDist_T_797; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_799 = fmt0_recA_rawIn_fractIn[312] ? 9'haf : _fmt0_recA_rawIn_normDist_T_798; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_800 = fmt0_recA_rawIn_fractIn[313] ? 9'hae : _fmt0_recA_rawIn_normDist_T_799; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_801 = fmt0_recA_rawIn_fractIn[314] ? 9'had : _fmt0_recA_rawIn_normDist_T_800; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_802 = fmt0_recA_rawIn_fractIn[315] ? 9'hac : _fmt0_recA_rawIn_normDist_T_801; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_803 = fmt0_recA_rawIn_fractIn[316] ? 9'hab : _fmt0_recA_rawIn_normDist_T_802; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_804 = fmt0_recA_rawIn_fractIn[317] ? 9'haa : _fmt0_recA_rawIn_normDist_T_803; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_805 = fmt0_recA_rawIn_fractIn[318] ? 9'ha9 : _fmt0_recA_rawIn_normDist_T_804; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_806 = fmt0_recA_rawIn_fractIn[319] ? 9'ha8 : _fmt0_recA_rawIn_normDist_T_805; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_807 = fmt0_recA_rawIn_fractIn[320] ? 9'ha7 : _fmt0_recA_rawIn_normDist_T_806; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_808 = fmt0_recA_rawIn_fractIn[321] ? 9'ha6 : _fmt0_recA_rawIn_normDist_T_807; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_809 = fmt0_recA_rawIn_fractIn[322] ? 9'ha5 : _fmt0_recA_rawIn_normDist_T_808; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_810 = fmt0_recA_rawIn_fractIn[323] ? 9'ha4 : _fmt0_recA_rawIn_normDist_T_809; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_811 = fmt0_recA_rawIn_fractIn[324] ? 9'ha3 : _fmt0_recA_rawIn_normDist_T_810; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_812 = fmt0_recA_rawIn_fractIn[325] ? 9'ha2 : _fmt0_recA_rawIn_normDist_T_811; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_813 = fmt0_recA_rawIn_fractIn[326] ? 9'ha1 : _fmt0_recA_rawIn_normDist_T_812; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_814 = fmt0_recA_rawIn_fractIn[327] ? 9'ha0 : _fmt0_recA_rawIn_normDist_T_813; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_815 = fmt0_recA_rawIn_fractIn[328] ? 9'h9f : _fmt0_recA_rawIn_normDist_T_814; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_816 = fmt0_recA_rawIn_fractIn[329] ? 9'h9e : _fmt0_recA_rawIn_normDist_T_815; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_817 = fmt0_recA_rawIn_fractIn[330] ? 9'h9d : _fmt0_recA_rawIn_normDist_T_816; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_818 = fmt0_recA_rawIn_fractIn[331] ? 9'h9c : _fmt0_recA_rawIn_normDist_T_817; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_819 = fmt0_recA_rawIn_fractIn[332] ? 9'h9b : _fmt0_recA_rawIn_normDist_T_818; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_820 = fmt0_recA_rawIn_fractIn[333] ? 9'h9a : _fmt0_recA_rawIn_normDist_T_819; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_821 = fmt0_recA_rawIn_fractIn[334] ? 9'h99 : _fmt0_recA_rawIn_normDist_T_820; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_822 = fmt0_recA_rawIn_fractIn[335] ? 9'h98 : _fmt0_recA_rawIn_normDist_T_821; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_823 = fmt0_recA_rawIn_fractIn[336] ? 9'h97 : _fmt0_recA_rawIn_normDist_T_822; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_824 = fmt0_recA_rawIn_fractIn[337] ? 9'h96 : _fmt0_recA_rawIn_normDist_T_823; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_825 = fmt0_recA_rawIn_fractIn[338] ? 9'h95 : _fmt0_recA_rawIn_normDist_T_824; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_826 = fmt0_recA_rawIn_fractIn[339] ? 9'h94 : _fmt0_recA_rawIn_normDist_T_825; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_827 = fmt0_recA_rawIn_fractIn[340] ? 9'h93 : _fmt0_recA_rawIn_normDist_T_826; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_828 = fmt0_recA_rawIn_fractIn[341] ? 9'h92 : _fmt0_recA_rawIn_normDist_T_827; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_829 = fmt0_recA_rawIn_fractIn[342] ? 9'h91 : _fmt0_recA_rawIn_normDist_T_828; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_830 = fmt0_recA_rawIn_fractIn[343] ? 9'h90 : _fmt0_recA_rawIn_normDist_T_829; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_831 = fmt0_recA_rawIn_fractIn[344] ? 9'h8f : _fmt0_recA_rawIn_normDist_T_830; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_832 = fmt0_recA_rawIn_fractIn[345] ? 9'h8e : _fmt0_recA_rawIn_normDist_T_831; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_833 = fmt0_recA_rawIn_fractIn[346] ? 9'h8d : _fmt0_recA_rawIn_normDist_T_832; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_834 = fmt0_recA_rawIn_fractIn[347] ? 9'h8c : _fmt0_recA_rawIn_normDist_T_833; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_835 = fmt0_recA_rawIn_fractIn[348] ? 9'h8b : _fmt0_recA_rawIn_normDist_T_834; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_836 = fmt0_recA_rawIn_fractIn[349] ? 9'h8a : _fmt0_recA_rawIn_normDist_T_835; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_837 = fmt0_recA_rawIn_fractIn[350] ? 9'h89 : _fmt0_recA_rawIn_normDist_T_836; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_838 = fmt0_recA_rawIn_fractIn[351] ? 9'h88 : _fmt0_recA_rawIn_normDist_T_837; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_839 = fmt0_recA_rawIn_fractIn[352] ? 9'h87 : _fmt0_recA_rawIn_normDist_T_838; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_840 = fmt0_recA_rawIn_fractIn[353] ? 9'h86 : _fmt0_recA_rawIn_normDist_T_839; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_841 = fmt0_recA_rawIn_fractIn[354] ? 9'h85 : _fmt0_recA_rawIn_normDist_T_840; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_842 = fmt0_recA_rawIn_fractIn[355] ? 9'h84 : _fmt0_recA_rawIn_normDist_T_841; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_843 = fmt0_recA_rawIn_fractIn[356] ? 9'h83 : _fmt0_recA_rawIn_normDist_T_842; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_844 = fmt0_recA_rawIn_fractIn[357] ? 9'h82 : _fmt0_recA_rawIn_normDist_T_843; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_845 = fmt0_recA_rawIn_fractIn[358] ? 9'h81 : _fmt0_recA_rawIn_normDist_T_844; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_846 = fmt0_recA_rawIn_fractIn[359] ? 9'h80 : _fmt0_recA_rawIn_normDist_T_845; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_847 = fmt0_recA_rawIn_fractIn[360] ? 9'h7f : _fmt0_recA_rawIn_normDist_T_846; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_848 = fmt0_recA_rawIn_fractIn[361] ? 9'h7e : _fmt0_recA_rawIn_normDist_T_847; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_849 = fmt0_recA_rawIn_fractIn[362] ? 9'h7d : _fmt0_recA_rawIn_normDist_T_848; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_850 = fmt0_recA_rawIn_fractIn[363] ? 9'h7c : _fmt0_recA_rawIn_normDist_T_849; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_851 = fmt0_recA_rawIn_fractIn[364] ? 9'h7b : _fmt0_recA_rawIn_normDist_T_850; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_852 = fmt0_recA_rawIn_fractIn[365] ? 9'h7a : _fmt0_recA_rawIn_normDist_T_851; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_853 = fmt0_recA_rawIn_fractIn[366] ? 9'h79 : _fmt0_recA_rawIn_normDist_T_852; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_854 = fmt0_recA_rawIn_fractIn[367] ? 9'h78 : _fmt0_recA_rawIn_normDist_T_853; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_855 = fmt0_recA_rawIn_fractIn[368] ? 9'h77 : _fmt0_recA_rawIn_normDist_T_854; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_856 = fmt0_recA_rawIn_fractIn[369] ? 9'h76 : _fmt0_recA_rawIn_normDist_T_855; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_857 = fmt0_recA_rawIn_fractIn[370] ? 9'h75 : _fmt0_recA_rawIn_normDist_T_856; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_858 = fmt0_recA_rawIn_fractIn[371] ? 9'h74 : _fmt0_recA_rawIn_normDist_T_857; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_859 = fmt0_recA_rawIn_fractIn[372] ? 9'h73 : _fmt0_recA_rawIn_normDist_T_858; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_860 = fmt0_recA_rawIn_fractIn[373] ? 9'h72 : _fmt0_recA_rawIn_normDist_T_859; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_861 = fmt0_recA_rawIn_fractIn[374] ? 9'h71 : _fmt0_recA_rawIn_normDist_T_860; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_862 = fmt0_recA_rawIn_fractIn[375] ? 9'h70 : _fmt0_recA_rawIn_normDist_T_861; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_863 = fmt0_recA_rawIn_fractIn[376] ? 9'h6f : _fmt0_recA_rawIn_normDist_T_862; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_864 = fmt0_recA_rawIn_fractIn[377] ? 9'h6e : _fmt0_recA_rawIn_normDist_T_863; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_865 = fmt0_recA_rawIn_fractIn[378] ? 9'h6d : _fmt0_recA_rawIn_normDist_T_864; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_866 = fmt0_recA_rawIn_fractIn[379] ? 9'h6c : _fmt0_recA_rawIn_normDist_T_865; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_867 = fmt0_recA_rawIn_fractIn[380] ? 9'h6b : _fmt0_recA_rawIn_normDist_T_866; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_868 = fmt0_recA_rawIn_fractIn[381] ? 9'h6a : _fmt0_recA_rawIn_normDist_T_867; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_869 = fmt0_recA_rawIn_fractIn[382] ? 9'h69 : _fmt0_recA_rawIn_normDist_T_868; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_870 = fmt0_recA_rawIn_fractIn[383] ? 9'h68 : _fmt0_recA_rawIn_normDist_T_869; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_871 = fmt0_recA_rawIn_fractIn[384] ? 9'h67 : _fmt0_recA_rawIn_normDist_T_870; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_872 = fmt0_recA_rawIn_fractIn[385] ? 9'h66 : _fmt0_recA_rawIn_normDist_T_871; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_873 = fmt0_recA_rawIn_fractIn[386] ? 9'h65 : _fmt0_recA_rawIn_normDist_T_872; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_874 = fmt0_recA_rawIn_fractIn[387] ? 9'h64 : _fmt0_recA_rawIn_normDist_T_873; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_875 = fmt0_recA_rawIn_fractIn[388] ? 9'h63 : _fmt0_recA_rawIn_normDist_T_874; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_876 = fmt0_recA_rawIn_fractIn[389] ? 9'h62 : _fmt0_recA_rawIn_normDist_T_875; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_877 = fmt0_recA_rawIn_fractIn[390] ? 9'h61 : _fmt0_recA_rawIn_normDist_T_876; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_878 = fmt0_recA_rawIn_fractIn[391] ? 9'h60 : _fmt0_recA_rawIn_normDist_T_877; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_879 = fmt0_recA_rawIn_fractIn[392] ? 9'h5f : _fmt0_recA_rawIn_normDist_T_878; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_880 = fmt0_recA_rawIn_fractIn[393] ? 9'h5e : _fmt0_recA_rawIn_normDist_T_879; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_881 = fmt0_recA_rawIn_fractIn[394] ? 9'h5d : _fmt0_recA_rawIn_normDist_T_880; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_882 = fmt0_recA_rawIn_fractIn[395] ? 9'h5c : _fmt0_recA_rawIn_normDist_T_881; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_883 = fmt0_recA_rawIn_fractIn[396] ? 9'h5b : _fmt0_recA_rawIn_normDist_T_882; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_884 = fmt0_recA_rawIn_fractIn[397] ? 9'h5a : _fmt0_recA_rawIn_normDist_T_883; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_885 = fmt0_recA_rawIn_fractIn[398] ? 9'h59 : _fmt0_recA_rawIn_normDist_T_884; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_886 = fmt0_recA_rawIn_fractIn[399] ? 9'h58 : _fmt0_recA_rawIn_normDist_T_885; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_887 = fmt0_recA_rawIn_fractIn[400] ? 9'h57 : _fmt0_recA_rawIn_normDist_T_886; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_888 = fmt0_recA_rawIn_fractIn[401] ? 9'h56 : _fmt0_recA_rawIn_normDist_T_887; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_889 = fmt0_recA_rawIn_fractIn[402] ? 9'h55 : _fmt0_recA_rawIn_normDist_T_888; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_890 = fmt0_recA_rawIn_fractIn[403] ? 9'h54 : _fmt0_recA_rawIn_normDist_T_889; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_891 = fmt0_recA_rawIn_fractIn[404] ? 9'h53 : _fmt0_recA_rawIn_normDist_T_890; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_892 = fmt0_recA_rawIn_fractIn[405] ? 9'h52 : _fmt0_recA_rawIn_normDist_T_891; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_893 = fmt0_recA_rawIn_fractIn[406] ? 9'h51 : _fmt0_recA_rawIn_normDist_T_892; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_894 = fmt0_recA_rawIn_fractIn[407] ? 9'h50 : _fmt0_recA_rawIn_normDist_T_893; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_895 = fmt0_recA_rawIn_fractIn[408] ? 9'h4f : _fmt0_recA_rawIn_normDist_T_894; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_896 = fmt0_recA_rawIn_fractIn[409] ? 9'h4e : _fmt0_recA_rawIn_normDist_T_895; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_897 = fmt0_recA_rawIn_fractIn[410] ? 9'h4d : _fmt0_recA_rawIn_normDist_T_896; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_898 = fmt0_recA_rawIn_fractIn[411] ? 9'h4c : _fmt0_recA_rawIn_normDist_T_897; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_899 = fmt0_recA_rawIn_fractIn[412] ? 9'h4b : _fmt0_recA_rawIn_normDist_T_898; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_900 = fmt0_recA_rawIn_fractIn[413] ? 9'h4a : _fmt0_recA_rawIn_normDist_T_899; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_901 = fmt0_recA_rawIn_fractIn[414] ? 9'h49 : _fmt0_recA_rawIn_normDist_T_900; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_902 = fmt0_recA_rawIn_fractIn[415] ? 9'h48 : _fmt0_recA_rawIn_normDist_T_901; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_903 = fmt0_recA_rawIn_fractIn[416] ? 9'h47 : _fmt0_recA_rawIn_normDist_T_902; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_904 = fmt0_recA_rawIn_fractIn[417] ? 9'h46 : _fmt0_recA_rawIn_normDist_T_903; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_905 = fmt0_recA_rawIn_fractIn[418] ? 9'h45 : _fmt0_recA_rawIn_normDist_T_904; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_906 = fmt0_recA_rawIn_fractIn[419] ? 9'h44 : _fmt0_recA_rawIn_normDist_T_905; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_907 = fmt0_recA_rawIn_fractIn[420] ? 9'h43 : _fmt0_recA_rawIn_normDist_T_906; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_908 = fmt0_recA_rawIn_fractIn[421] ? 9'h42 : _fmt0_recA_rawIn_normDist_T_907; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_909 = fmt0_recA_rawIn_fractIn[422] ? 9'h41 : _fmt0_recA_rawIn_normDist_T_908; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_910 = fmt0_recA_rawIn_fractIn[423] ? 9'h40 : _fmt0_recA_rawIn_normDist_T_909; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_911 = fmt0_recA_rawIn_fractIn[424] ? 9'h3f : _fmt0_recA_rawIn_normDist_T_910; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_912 = fmt0_recA_rawIn_fractIn[425] ? 9'h3e : _fmt0_recA_rawIn_normDist_T_911; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_913 = fmt0_recA_rawIn_fractIn[426] ? 9'h3d : _fmt0_recA_rawIn_normDist_T_912; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_914 = fmt0_recA_rawIn_fractIn[427] ? 9'h3c : _fmt0_recA_rawIn_normDist_T_913; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_915 = fmt0_recA_rawIn_fractIn[428] ? 9'h3b : _fmt0_recA_rawIn_normDist_T_914; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_916 = fmt0_recA_rawIn_fractIn[429] ? 9'h3a : _fmt0_recA_rawIn_normDist_T_915; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_917 = fmt0_recA_rawIn_fractIn[430] ? 9'h39 : _fmt0_recA_rawIn_normDist_T_916; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_918 = fmt0_recA_rawIn_fractIn[431] ? 9'h38 : _fmt0_recA_rawIn_normDist_T_917; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_919 = fmt0_recA_rawIn_fractIn[432] ? 9'h37 : _fmt0_recA_rawIn_normDist_T_918; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_920 = fmt0_recA_rawIn_fractIn[433] ? 9'h36 : _fmt0_recA_rawIn_normDist_T_919; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_921 = fmt0_recA_rawIn_fractIn[434] ? 9'h35 : _fmt0_recA_rawIn_normDist_T_920; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_922 = fmt0_recA_rawIn_fractIn[435] ? 9'h34 : _fmt0_recA_rawIn_normDist_T_921; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_923 = fmt0_recA_rawIn_fractIn[436] ? 9'h33 : _fmt0_recA_rawIn_normDist_T_922; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_924 = fmt0_recA_rawIn_fractIn[437] ? 9'h32 : _fmt0_recA_rawIn_normDist_T_923; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_925 = fmt0_recA_rawIn_fractIn[438] ? 9'h31 : _fmt0_recA_rawIn_normDist_T_924; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_926 = fmt0_recA_rawIn_fractIn[439] ? 9'h30 : _fmt0_recA_rawIn_normDist_T_925; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_927 = fmt0_recA_rawIn_fractIn[440] ? 9'h2f : _fmt0_recA_rawIn_normDist_T_926; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_928 = fmt0_recA_rawIn_fractIn[441] ? 9'h2e : _fmt0_recA_rawIn_normDist_T_927; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_929 = fmt0_recA_rawIn_fractIn[442] ? 9'h2d : _fmt0_recA_rawIn_normDist_T_928; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_930 = fmt0_recA_rawIn_fractIn[443] ? 9'h2c : _fmt0_recA_rawIn_normDist_T_929; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_931 = fmt0_recA_rawIn_fractIn[444] ? 9'h2b : _fmt0_recA_rawIn_normDist_T_930; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_932 = fmt0_recA_rawIn_fractIn[445] ? 9'h2a : _fmt0_recA_rawIn_normDist_T_931; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_933 = fmt0_recA_rawIn_fractIn[446] ? 9'h29 : _fmt0_recA_rawIn_normDist_T_932; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_934 = fmt0_recA_rawIn_fractIn[447] ? 9'h28 : _fmt0_recA_rawIn_normDist_T_933; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_935 = fmt0_recA_rawIn_fractIn[448] ? 9'h27 : _fmt0_recA_rawIn_normDist_T_934; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_936 = fmt0_recA_rawIn_fractIn[449] ? 9'h26 : _fmt0_recA_rawIn_normDist_T_935; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_937 = fmt0_recA_rawIn_fractIn[450] ? 9'h25 : _fmt0_recA_rawIn_normDist_T_936; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_938 = fmt0_recA_rawIn_fractIn[451] ? 9'h24 : _fmt0_recA_rawIn_normDist_T_937; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_939 = fmt0_recA_rawIn_fractIn[452] ? 9'h23 : _fmt0_recA_rawIn_normDist_T_938; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_940 = fmt0_recA_rawIn_fractIn[453] ? 9'h22 : _fmt0_recA_rawIn_normDist_T_939; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_941 = fmt0_recA_rawIn_fractIn[454] ? 9'h21 : _fmt0_recA_rawIn_normDist_T_940; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_942 = fmt0_recA_rawIn_fractIn[455] ? 9'h20 : _fmt0_recA_rawIn_normDist_T_941; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_943 = fmt0_recA_rawIn_fractIn[456] ? 9'h1f : _fmt0_recA_rawIn_normDist_T_942; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_944 = fmt0_recA_rawIn_fractIn[457] ? 9'h1e : _fmt0_recA_rawIn_normDist_T_943; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_945 = fmt0_recA_rawIn_fractIn[458] ? 9'h1d : _fmt0_recA_rawIn_normDist_T_944; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_946 = fmt0_recA_rawIn_fractIn[459] ? 9'h1c : _fmt0_recA_rawIn_normDist_T_945; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_947 = fmt0_recA_rawIn_fractIn[460] ? 9'h1b : _fmt0_recA_rawIn_normDist_T_946; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_948 = fmt0_recA_rawIn_fractIn[461] ? 9'h1a : _fmt0_recA_rawIn_normDist_T_947; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_949 = fmt0_recA_rawIn_fractIn[462] ? 9'h19 : _fmt0_recA_rawIn_normDist_T_948; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_950 = fmt0_recA_rawIn_fractIn[463] ? 9'h18 : _fmt0_recA_rawIn_normDist_T_949; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_951 = fmt0_recA_rawIn_fractIn[464] ? 9'h17 : _fmt0_recA_rawIn_normDist_T_950; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_952 = fmt0_recA_rawIn_fractIn[465] ? 9'h16 : _fmt0_recA_rawIn_normDist_T_951; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_953 = fmt0_recA_rawIn_fractIn[466] ? 9'h15 : _fmt0_recA_rawIn_normDist_T_952; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_954 = fmt0_recA_rawIn_fractIn[467] ? 9'h14 : _fmt0_recA_rawIn_normDist_T_953; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_955 = fmt0_recA_rawIn_fractIn[468] ? 9'h13 : _fmt0_recA_rawIn_normDist_T_954; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_956 = fmt0_recA_rawIn_fractIn[469] ? 9'h12 : _fmt0_recA_rawIn_normDist_T_955; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_957 = fmt0_recA_rawIn_fractIn[470] ? 9'h11 : _fmt0_recA_rawIn_normDist_T_956; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_958 = fmt0_recA_rawIn_fractIn[471] ? 9'h10 : _fmt0_recA_rawIn_normDist_T_957; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_959 = fmt0_recA_rawIn_fractIn[472] ? 9'hf : _fmt0_recA_rawIn_normDist_T_958; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_960 = fmt0_recA_rawIn_fractIn[473] ? 9'he : _fmt0_recA_rawIn_normDist_T_959; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_961 = fmt0_recA_rawIn_fractIn[474] ? 9'hd : _fmt0_recA_rawIn_normDist_T_960; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_962 = fmt0_recA_rawIn_fractIn[475] ? 9'hc : _fmt0_recA_rawIn_normDist_T_961; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_963 = fmt0_recA_rawIn_fractIn[476] ? 9'hb : _fmt0_recA_rawIn_normDist_T_962; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_964 = fmt0_recA_rawIn_fractIn[477] ? 9'ha : _fmt0_recA_rawIn_normDist_T_963; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_965 = fmt0_recA_rawIn_fractIn[478] ? 9'h9 : _fmt0_recA_rawIn_normDist_T_964; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_966 = fmt0_recA_rawIn_fractIn[479] ? 9'h8 : _fmt0_recA_rawIn_normDist_T_965; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_967 = fmt0_recA_rawIn_fractIn[480] ? 9'h7 : _fmt0_recA_rawIn_normDist_T_966; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_968 = fmt0_recA_rawIn_fractIn[481] ? 9'h6 : _fmt0_recA_rawIn_normDist_T_967; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_969 = fmt0_recA_rawIn_fractIn[482] ? 9'h5 : _fmt0_recA_rawIn_normDist_T_968; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_970 = fmt0_recA_rawIn_fractIn[483] ? 9'h4 : _fmt0_recA_rawIn_normDist_T_969; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_971 = fmt0_recA_rawIn_fractIn[484] ? 9'h3 : _fmt0_recA_rawIn_normDist_T_970; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_972 = fmt0_recA_rawIn_fractIn[485] ? 9'h2 : _fmt0_recA_rawIn_normDist_T_971; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recA_rawIn_normDist_T_973 = fmt0_recA_rawIn_fractIn[486] ? 9'h1 : _fmt0_recA_rawIn_normDist_T_972; // @[Mux.scala 47:70]
  wire [8:0] fmt0_recA_rawIn_normDist = fmt0_recA_rawIn_fractIn[487] ? 9'h0 : _fmt0_recA_rawIn_normDist_T_973; // @[Mux.scala 47:70]
  wire [998:0] _GEN_4 = {{511'd0}, fmt0_recA_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [998:0] _fmt0_recA_rawIn_subnormFract_T = _GEN_4 << fmt0_recA_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [487:0] fmt0_recA_rawIn_subnormFract = {_fmt0_recA_rawIn_subnormFract_T[486:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [23:0] _GEN_9 = {{15'd0}, fmt0_recA_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [23:0] _fmt0_recA_rawIn_adjustedExp_T = _GEN_9 ^ 24'hffffff; // @[rawFloatFromFN.scala 55:18]
  wire [23:0] _fmt0_recA_rawIn_adjustedExp_T_1 = fmt0_recA_rawIn_isZeroExpIn ? _fmt0_recA_rawIn_adjustedExp_T : {{1
    'd0}, fmt0_recA_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _fmt0_recA_rawIn_adjustedExp_T_2 = fmt0_recA_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [22:0] _GEN_10 = {{21'd0}, _fmt0_recA_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [22:0] _fmt0_recA_rawIn_adjustedExp_T_3 = 23'h400000 | _GEN_10; // @[rawFloatFromFN.scala 58:9]
  wire [23:0] _GEN_11 = {{1'd0}, _fmt0_recA_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [23:0] fmt0_recA_rawIn_adjustedExp = _fmt0_recA_rawIn_adjustedExp_T_1 + _GEN_11; // @[rawFloatFromFN.scala 57:9]
  wire  fmt0_recA_rawIn_isZero = fmt0_recA_rawIn_isZeroExpIn & fmt0_recA_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  fmt0_recA_rawIn_isSpecial = fmt0_recA_rawIn_adjustedExp[23:22] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  fmt0_recA_rawIn__isNaN = fmt0_recA_rawIn_isSpecial & ~fmt0_recA_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [24:0] fmt0_recA_rawIn__sExp = {1'b0,$signed(fmt0_recA_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _fmt0_recA_rawIn_out_sig_T = ~fmt0_recA_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [487:0] _fmt0_recA_rawIn_out_sig_T_2 = fmt0_recA_rawIn_isZeroExpIn ? fmt0_recA_rawIn_subnormFract :
    fmt0_recA_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [489:0] fmt0_recA_rawIn__sig = {1'h0,_fmt0_recA_rawIn_out_sig_T,_fmt0_recA_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _fmt0_recA_T_2 = fmt0_recA_rawIn_isZero ? 3'h0 : fmt0_recA_rawIn__sExp[23:21]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_12 = {{2'd0}, fmt0_recA_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _fmt0_recA_T_4 = _fmt0_recA_T_2 | _GEN_12; // @[recFNFromFN.scala 48:76]
  wire [24:0] _fmt0_recA_T_7 = {fmt0_recA_rawIn_sign,_fmt0_recA_T_4,fmt0_recA_rawIn__sExp[20:0]}; // @[recFNFromFN.scala 49:45]
  wire  fmt0_recB_rawIn_sign = io_b[511]; // @[rawFloatFromFN.scala 44:18]
  wire [22:0] fmt0_recB_rawIn_expIn = io_b[510:488]; // @[rawFloatFromFN.scala 45:19]
  wire [487:0] fmt0_recB_rawIn_fractIn = io_b[487:0]; // @[rawFloatFromFN.scala 46:21]
  wire  fmt0_recB_rawIn_isZeroExpIn = fmt0_recB_rawIn_expIn == 23'h0; // @[rawFloatFromFN.scala 48:30]
  wire  fmt0_recB_rawIn_isZeroFractIn = fmt0_recB_rawIn_fractIn == 488'h0; // @[rawFloatFromFN.scala 49:34]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_488 = fmt0_recB_rawIn_fractIn[1] ? 9'h1e6 : 9'h1e7; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_489 = fmt0_recB_rawIn_fractIn[2] ? 9'h1e5 : _fmt0_recB_rawIn_normDist_T_488; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_490 = fmt0_recB_rawIn_fractIn[3] ? 9'h1e4 : _fmt0_recB_rawIn_normDist_T_489; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_491 = fmt0_recB_rawIn_fractIn[4] ? 9'h1e3 : _fmt0_recB_rawIn_normDist_T_490; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_492 = fmt0_recB_rawIn_fractIn[5] ? 9'h1e2 : _fmt0_recB_rawIn_normDist_T_491; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_493 = fmt0_recB_rawIn_fractIn[6] ? 9'h1e1 : _fmt0_recB_rawIn_normDist_T_492; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_494 = fmt0_recB_rawIn_fractIn[7] ? 9'h1e0 : _fmt0_recB_rawIn_normDist_T_493; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_495 = fmt0_recB_rawIn_fractIn[8] ? 9'h1df : _fmt0_recB_rawIn_normDist_T_494; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_496 = fmt0_recB_rawIn_fractIn[9] ? 9'h1de : _fmt0_recB_rawIn_normDist_T_495; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_497 = fmt0_recB_rawIn_fractIn[10] ? 9'h1dd : _fmt0_recB_rawIn_normDist_T_496; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_498 = fmt0_recB_rawIn_fractIn[11] ? 9'h1dc : _fmt0_recB_rawIn_normDist_T_497; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_499 = fmt0_recB_rawIn_fractIn[12] ? 9'h1db : _fmt0_recB_rawIn_normDist_T_498; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_500 = fmt0_recB_rawIn_fractIn[13] ? 9'h1da : _fmt0_recB_rawIn_normDist_T_499; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_501 = fmt0_recB_rawIn_fractIn[14] ? 9'h1d9 : _fmt0_recB_rawIn_normDist_T_500; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_502 = fmt0_recB_rawIn_fractIn[15] ? 9'h1d8 : _fmt0_recB_rawIn_normDist_T_501; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_503 = fmt0_recB_rawIn_fractIn[16] ? 9'h1d7 : _fmt0_recB_rawIn_normDist_T_502; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_504 = fmt0_recB_rawIn_fractIn[17] ? 9'h1d6 : _fmt0_recB_rawIn_normDist_T_503; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_505 = fmt0_recB_rawIn_fractIn[18] ? 9'h1d5 : _fmt0_recB_rawIn_normDist_T_504; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_506 = fmt0_recB_rawIn_fractIn[19] ? 9'h1d4 : _fmt0_recB_rawIn_normDist_T_505; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_507 = fmt0_recB_rawIn_fractIn[20] ? 9'h1d3 : _fmt0_recB_rawIn_normDist_T_506; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_508 = fmt0_recB_rawIn_fractIn[21] ? 9'h1d2 : _fmt0_recB_rawIn_normDist_T_507; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_509 = fmt0_recB_rawIn_fractIn[22] ? 9'h1d1 : _fmt0_recB_rawIn_normDist_T_508; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_510 = fmt0_recB_rawIn_fractIn[23] ? 9'h1d0 : _fmt0_recB_rawIn_normDist_T_509; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_511 = fmt0_recB_rawIn_fractIn[24] ? 9'h1cf : _fmt0_recB_rawIn_normDist_T_510; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_512 = fmt0_recB_rawIn_fractIn[25] ? 9'h1ce : _fmt0_recB_rawIn_normDist_T_511; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_513 = fmt0_recB_rawIn_fractIn[26] ? 9'h1cd : _fmt0_recB_rawIn_normDist_T_512; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_514 = fmt0_recB_rawIn_fractIn[27] ? 9'h1cc : _fmt0_recB_rawIn_normDist_T_513; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_515 = fmt0_recB_rawIn_fractIn[28] ? 9'h1cb : _fmt0_recB_rawIn_normDist_T_514; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_516 = fmt0_recB_rawIn_fractIn[29] ? 9'h1ca : _fmt0_recB_rawIn_normDist_T_515; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_517 = fmt0_recB_rawIn_fractIn[30] ? 9'h1c9 : _fmt0_recB_rawIn_normDist_T_516; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_518 = fmt0_recB_rawIn_fractIn[31] ? 9'h1c8 : _fmt0_recB_rawIn_normDist_T_517; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_519 = fmt0_recB_rawIn_fractIn[32] ? 9'h1c7 : _fmt0_recB_rawIn_normDist_T_518; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_520 = fmt0_recB_rawIn_fractIn[33] ? 9'h1c6 : _fmt0_recB_rawIn_normDist_T_519; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_521 = fmt0_recB_rawIn_fractIn[34] ? 9'h1c5 : _fmt0_recB_rawIn_normDist_T_520; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_522 = fmt0_recB_rawIn_fractIn[35] ? 9'h1c4 : _fmt0_recB_rawIn_normDist_T_521; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_523 = fmt0_recB_rawIn_fractIn[36] ? 9'h1c3 : _fmt0_recB_rawIn_normDist_T_522; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_524 = fmt0_recB_rawIn_fractIn[37] ? 9'h1c2 : _fmt0_recB_rawIn_normDist_T_523; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_525 = fmt0_recB_rawIn_fractIn[38] ? 9'h1c1 : _fmt0_recB_rawIn_normDist_T_524; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_526 = fmt0_recB_rawIn_fractIn[39] ? 9'h1c0 : _fmt0_recB_rawIn_normDist_T_525; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_527 = fmt0_recB_rawIn_fractIn[40] ? 9'h1bf : _fmt0_recB_rawIn_normDist_T_526; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_528 = fmt0_recB_rawIn_fractIn[41] ? 9'h1be : _fmt0_recB_rawIn_normDist_T_527; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_529 = fmt0_recB_rawIn_fractIn[42] ? 9'h1bd : _fmt0_recB_rawIn_normDist_T_528; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_530 = fmt0_recB_rawIn_fractIn[43] ? 9'h1bc : _fmt0_recB_rawIn_normDist_T_529; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_531 = fmt0_recB_rawIn_fractIn[44] ? 9'h1bb : _fmt0_recB_rawIn_normDist_T_530; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_532 = fmt0_recB_rawIn_fractIn[45] ? 9'h1ba : _fmt0_recB_rawIn_normDist_T_531; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_533 = fmt0_recB_rawIn_fractIn[46] ? 9'h1b9 : _fmt0_recB_rawIn_normDist_T_532; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_534 = fmt0_recB_rawIn_fractIn[47] ? 9'h1b8 : _fmt0_recB_rawIn_normDist_T_533; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_535 = fmt0_recB_rawIn_fractIn[48] ? 9'h1b7 : _fmt0_recB_rawIn_normDist_T_534; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_536 = fmt0_recB_rawIn_fractIn[49] ? 9'h1b6 : _fmt0_recB_rawIn_normDist_T_535; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_537 = fmt0_recB_rawIn_fractIn[50] ? 9'h1b5 : _fmt0_recB_rawIn_normDist_T_536; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_538 = fmt0_recB_rawIn_fractIn[51] ? 9'h1b4 : _fmt0_recB_rawIn_normDist_T_537; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_539 = fmt0_recB_rawIn_fractIn[52] ? 9'h1b3 : _fmt0_recB_rawIn_normDist_T_538; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_540 = fmt0_recB_rawIn_fractIn[53] ? 9'h1b2 : _fmt0_recB_rawIn_normDist_T_539; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_541 = fmt0_recB_rawIn_fractIn[54] ? 9'h1b1 : _fmt0_recB_rawIn_normDist_T_540; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_542 = fmt0_recB_rawIn_fractIn[55] ? 9'h1b0 : _fmt0_recB_rawIn_normDist_T_541; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_543 = fmt0_recB_rawIn_fractIn[56] ? 9'h1af : _fmt0_recB_rawIn_normDist_T_542; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_544 = fmt0_recB_rawIn_fractIn[57] ? 9'h1ae : _fmt0_recB_rawIn_normDist_T_543; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_545 = fmt0_recB_rawIn_fractIn[58] ? 9'h1ad : _fmt0_recB_rawIn_normDist_T_544; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_546 = fmt0_recB_rawIn_fractIn[59] ? 9'h1ac : _fmt0_recB_rawIn_normDist_T_545; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_547 = fmt0_recB_rawIn_fractIn[60] ? 9'h1ab : _fmt0_recB_rawIn_normDist_T_546; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_548 = fmt0_recB_rawIn_fractIn[61] ? 9'h1aa : _fmt0_recB_rawIn_normDist_T_547; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_549 = fmt0_recB_rawIn_fractIn[62] ? 9'h1a9 : _fmt0_recB_rawIn_normDist_T_548; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_550 = fmt0_recB_rawIn_fractIn[63] ? 9'h1a8 : _fmt0_recB_rawIn_normDist_T_549; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_551 = fmt0_recB_rawIn_fractIn[64] ? 9'h1a7 : _fmt0_recB_rawIn_normDist_T_550; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_552 = fmt0_recB_rawIn_fractIn[65] ? 9'h1a6 : _fmt0_recB_rawIn_normDist_T_551; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_553 = fmt0_recB_rawIn_fractIn[66] ? 9'h1a5 : _fmt0_recB_rawIn_normDist_T_552; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_554 = fmt0_recB_rawIn_fractIn[67] ? 9'h1a4 : _fmt0_recB_rawIn_normDist_T_553; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_555 = fmt0_recB_rawIn_fractIn[68] ? 9'h1a3 : _fmt0_recB_rawIn_normDist_T_554; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_556 = fmt0_recB_rawIn_fractIn[69] ? 9'h1a2 : _fmt0_recB_rawIn_normDist_T_555; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_557 = fmt0_recB_rawIn_fractIn[70] ? 9'h1a1 : _fmt0_recB_rawIn_normDist_T_556; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_558 = fmt0_recB_rawIn_fractIn[71] ? 9'h1a0 : _fmt0_recB_rawIn_normDist_T_557; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_559 = fmt0_recB_rawIn_fractIn[72] ? 9'h19f : _fmt0_recB_rawIn_normDist_T_558; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_560 = fmt0_recB_rawIn_fractIn[73] ? 9'h19e : _fmt0_recB_rawIn_normDist_T_559; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_561 = fmt0_recB_rawIn_fractIn[74] ? 9'h19d : _fmt0_recB_rawIn_normDist_T_560; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_562 = fmt0_recB_rawIn_fractIn[75] ? 9'h19c : _fmt0_recB_rawIn_normDist_T_561; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_563 = fmt0_recB_rawIn_fractIn[76] ? 9'h19b : _fmt0_recB_rawIn_normDist_T_562; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_564 = fmt0_recB_rawIn_fractIn[77] ? 9'h19a : _fmt0_recB_rawIn_normDist_T_563; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_565 = fmt0_recB_rawIn_fractIn[78] ? 9'h199 : _fmt0_recB_rawIn_normDist_T_564; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_566 = fmt0_recB_rawIn_fractIn[79] ? 9'h198 : _fmt0_recB_rawIn_normDist_T_565; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_567 = fmt0_recB_rawIn_fractIn[80] ? 9'h197 : _fmt0_recB_rawIn_normDist_T_566; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_568 = fmt0_recB_rawIn_fractIn[81] ? 9'h196 : _fmt0_recB_rawIn_normDist_T_567; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_569 = fmt0_recB_rawIn_fractIn[82] ? 9'h195 : _fmt0_recB_rawIn_normDist_T_568; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_570 = fmt0_recB_rawIn_fractIn[83] ? 9'h194 : _fmt0_recB_rawIn_normDist_T_569; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_571 = fmt0_recB_rawIn_fractIn[84] ? 9'h193 : _fmt0_recB_rawIn_normDist_T_570; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_572 = fmt0_recB_rawIn_fractIn[85] ? 9'h192 : _fmt0_recB_rawIn_normDist_T_571; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_573 = fmt0_recB_rawIn_fractIn[86] ? 9'h191 : _fmt0_recB_rawIn_normDist_T_572; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_574 = fmt0_recB_rawIn_fractIn[87] ? 9'h190 : _fmt0_recB_rawIn_normDist_T_573; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_575 = fmt0_recB_rawIn_fractIn[88] ? 9'h18f : _fmt0_recB_rawIn_normDist_T_574; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_576 = fmt0_recB_rawIn_fractIn[89] ? 9'h18e : _fmt0_recB_rawIn_normDist_T_575; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_577 = fmt0_recB_rawIn_fractIn[90] ? 9'h18d : _fmt0_recB_rawIn_normDist_T_576; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_578 = fmt0_recB_rawIn_fractIn[91] ? 9'h18c : _fmt0_recB_rawIn_normDist_T_577; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_579 = fmt0_recB_rawIn_fractIn[92] ? 9'h18b : _fmt0_recB_rawIn_normDist_T_578; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_580 = fmt0_recB_rawIn_fractIn[93] ? 9'h18a : _fmt0_recB_rawIn_normDist_T_579; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_581 = fmt0_recB_rawIn_fractIn[94] ? 9'h189 : _fmt0_recB_rawIn_normDist_T_580; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_582 = fmt0_recB_rawIn_fractIn[95] ? 9'h188 : _fmt0_recB_rawIn_normDist_T_581; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_583 = fmt0_recB_rawIn_fractIn[96] ? 9'h187 : _fmt0_recB_rawIn_normDist_T_582; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_584 = fmt0_recB_rawIn_fractIn[97] ? 9'h186 : _fmt0_recB_rawIn_normDist_T_583; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_585 = fmt0_recB_rawIn_fractIn[98] ? 9'h185 : _fmt0_recB_rawIn_normDist_T_584; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_586 = fmt0_recB_rawIn_fractIn[99] ? 9'h184 : _fmt0_recB_rawIn_normDist_T_585; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_587 = fmt0_recB_rawIn_fractIn[100] ? 9'h183 : _fmt0_recB_rawIn_normDist_T_586; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_588 = fmt0_recB_rawIn_fractIn[101] ? 9'h182 : _fmt0_recB_rawIn_normDist_T_587; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_589 = fmt0_recB_rawIn_fractIn[102] ? 9'h181 : _fmt0_recB_rawIn_normDist_T_588; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_590 = fmt0_recB_rawIn_fractIn[103] ? 9'h180 : _fmt0_recB_rawIn_normDist_T_589; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_591 = fmt0_recB_rawIn_fractIn[104] ? 9'h17f : _fmt0_recB_rawIn_normDist_T_590; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_592 = fmt0_recB_rawIn_fractIn[105] ? 9'h17e : _fmt0_recB_rawIn_normDist_T_591; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_593 = fmt0_recB_rawIn_fractIn[106] ? 9'h17d : _fmt0_recB_rawIn_normDist_T_592; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_594 = fmt0_recB_rawIn_fractIn[107] ? 9'h17c : _fmt0_recB_rawIn_normDist_T_593; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_595 = fmt0_recB_rawIn_fractIn[108] ? 9'h17b : _fmt0_recB_rawIn_normDist_T_594; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_596 = fmt0_recB_rawIn_fractIn[109] ? 9'h17a : _fmt0_recB_rawIn_normDist_T_595; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_597 = fmt0_recB_rawIn_fractIn[110] ? 9'h179 : _fmt0_recB_rawIn_normDist_T_596; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_598 = fmt0_recB_rawIn_fractIn[111] ? 9'h178 : _fmt0_recB_rawIn_normDist_T_597; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_599 = fmt0_recB_rawIn_fractIn[112] ? 9'h177 : _fmt0_recB_rawIn_normDist_T_598; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_600 = fmt0_recB_rawIn_fractIn[113] ? 9'h176 : _fmt0_recB_rawIn_normDist_T_599; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_601 = fmt0_recB_rawIn_fractIn[114] ? 9'h175 : _fmt0_recB_rawIn_normDist_T_600; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_602 = fmt0_recB_rawIn_fractIn[115] ? 9'h174 : _fmt0_recB_rawIn_normDist_T_601; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_603 = fmt0_recB_rawIn_fractIn[116] ? 9'h173 : _fmt0_recB_rawIn_normDist_T_602; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_604 = fmt0_recB_rawIn_fractIn[117] ? 9'h172 : _fmt0_recB_rawIn_normDist_T_603; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_605 = fmt0_recB_rawIn_fractIn[118] ? 9'h171 : _fmt0_recB_rawIn_normDist_T_604; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_606 = fmt0_recB_rawIn_fractIn[119] ? 9'h170 : _fmt0_recB_rawIn_normDist_T_605; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_607 = fmt0_recB_rawIn_fractIn[120] ? 9'h16f : _fmt0_recB_rawIn_normDist_T_606; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_608 = fmt0_recB_rawIn_fractIn[121] ? 9'h16e : _fmt0_recB_rawIn_normDist_T_607; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_609 = fmt0_recB_rawIn_fractIn[122] ? 9'h16d : _fmt0_recB_rawIn_normDist_T_608; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_610 = fmt0_recB_rawIn_fractIn[123] ? 9'h16c : _fmt0_recB_rawIn_normDist_T_609; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_611 = fmt0_recB_rawIn_fractIn[124] ? 9'h16b : _fmt0_recB_rawIn_normDist_T_610; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_612 = fmt0_recB_rawIn_fractIn[125] ? 9'h16a : _fmt0_recB_rawIn_normDist_T_611; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_613 = fmt0_recB_rawIn_fractIn[126] ? 9'h169 : _fmt0_recB_rawIn_normDist_T_612; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_614 = fmt0_recB_rawIn_fractIn[127] ? 9'h168 : _fmt0_recB_rawIn_normDist_T_613; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_615 = fmt0_recB_rawIn_fractIn[128] ? 9'h167 : _fmt0_recB_rawIn_normDist_T_614; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_616 = fmt0_recB_rawIn_fractIn[129] ? 9'h166 : _fmt0_recB_rawIn_normDist_T_615; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_617 = fmt0_recB_rawIn_fractIn[130] ? 9'h165 : _fmt0_recB_rawIn_normDist_T_616; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_618 = fmt0_recB_rawIn_fractIn[131] ? 9'h164 : _fmt0_recB_rawIn_normDist_T_617; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_619 = fmt0_recB_rawIn_fractIn[132] ? 9'h163 : _fmt0_recB_rawIn_normDist_T_618; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_620 = fmt0_recB_rawIn_fractIn[133] ? 9'h162 : _fmt0_recB_rawIn_normDist_T_619; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_621 = fmt0_recB_rawIn_fractIn[134] ? 9'h161 : _fmt0_recB_rawIn_normDist_T_620; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_622 = fmt0_recB_rawIn_fractIn[135] ? 9'h160 : _fmt0_recB_rawIn_normDist_T_621; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_623 = fmt0_recB_rawIn_fractIn[136] ? 9'h15f : _fmt0_recB_rawIn_normDist_T_622; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_624 = fmt0_recB_rawIn_fractIn[137] ? 9'h15e : _fmt0_recB_rawIn_normDist_T_623; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_625 = fmt0_recB_rawIn_fractIn[138] ? 9'h15d : _fmt0_recB_rawIn_normDist_T_624; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_626 = fmt0_recB_rawIn_fractIn[139] ? 9'h15c : _fmt0_recB_rawIn_normDist_T_625; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_627 = fmt0_recB_rawIn_fractIn[140] ? 9'h15b : _fmt0_recB_rawIn_normDist_T_626; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_628 = fmt0_recB_rawIn_fractIn[141] ? 9'h15a : _fmt0_recB_rawIn_normDist_T_627; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_629 = fmt0_recB_rawIn_fractIn[142] ? 9'h159 : _fmt0_recB_rawIn_normDist_T_628; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_630 = fmt0_recB_rawIn_fractIn[143] ? 9'h158 : _fmt0_recB_rawIn_normDist_T_629; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_631 = fmt0_recB_rawIn_fractIn[144] ? 9'h157 : _fmt0_recB_rawIn_normDist_T_630; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_632 = fmt0_recB_rawIn_fractIn[145] ? 9'h156 : _fmt0_recB_rawIn_normDist_T_631; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_633 = fmt0_recB_rawIn_fractIn[146] ? 9'h155 : _fmt0_recB_rawIn_normDist_T_632; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_634 = fmt0_recB_rawIn_fractIn[147] ? 9'h154 : _fmt0_recB_rawIn_normDist_T_633; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_635 = fmt0_recB_rawIn_fractIn[148] ? 9'h153 : _fmt0_recB_rawIn_normDist_T_634; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_636 = fmt0_recB_rawIn_fractIn[149] ? 9'h152 : _fmt0_recB_rawIn_normDist_T_635; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_637 = fmt0_recB_rawIn_fractIn[150] ? 9'h151 : _fmt0_recB_rawIn_normDist_T_636; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_638 = fmt0_recB_rawIn_fractIn[151] ? 9'h150 : _fmt0_recB_rawIn_normDist_T_637; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_639 = fmt0_recB_rawIn_fractIn[152] ? 9'h14f : _fmt0_recB_rawIn_normDist_T_638; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_640 = fmt0_recB_rawIn_fractIn[153] ? 9'h14e : _fmt0_recB_rawIn_normDist_T_639; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_641 = fmt0_recB_rawIn_fractIn[154] ? 9'h14d : _fmt0_recB_rawIn_normDist_T_640; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_642 = fmt0_recB_rawIn_fractIn[155] ? 9'h14c : _fmt0_recB_rawIn_normDist_T_641; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_643 = fmt0_recB_rawIn_fractIn[156] ? 9'h14b : _fmt0_recB_rawIn_normDist_T_642; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_644 = fmt0_recB_rawIn_fractIn[157] ? 9'h14a : _fmt0_recB_rawIn_normDist_T_643; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_645 = fmt0_recB_rawIn_fractIn[158] ? 9'h149 : _fmt0_recB_rawIn_normDist_T_644; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_646 = fmt0_recB_rawIn_fractIn[159] ? 9'h148 : _fmt0_recB_rawIn_normDist_T_645; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_647 = fmt0_recB_rawIn_fractIn[160] ? 9'h147 : _fmt0_recB_rawIn_normDist_T_646; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_648 = fmt0_recB_rawIn_fractIn[161] ? 9'h146 : _fmt0_recB_rawIn_normDist_T_647; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_649 = fmt0_recB_rawIn_fractIn[162] ? 9'h145 : _fmt0_recB_rawIn_normDist_T_648; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_650 = fmt0_recB_rawIn_fractIn[163] ? 9'h144 : _fmt0_recB_rawIn_normDist_T_649; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_651 = fmt0_recB_rawIn_fractIn[164] ? 9'h143 : _fmt0_recB_rawIn_normDist_T_650; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_652 = fmt0_recB_rawIn_fractIn[165] ? 9'h142 : _fmt0_recB_rawIn_normDist_T_651; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_653 = fmt0_recB_rawIn_fractIn[166] ? 9'h141 : _fmt0_recB_rawIn_normDist_T_652; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_654 = fmt0_recB_rawIn_fractIn[167] ? 9'h140 : _fmt0_recB_rawIn_normDist_T_653; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_655 = fmt0_recB_rawIn_fractIn[168] ? 9'h13f : _fmt0_recB_rawIn_normDist_T_654; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_656 = fmt0_recB_rawIn_fractIn[169] ? 9'h13e : _fmt0_recB_rawIn_normDist_T_655; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_657 = fmt0_recB_rawIn_fractIn[170] ? 9'h13d : _fmt0_recB_rawIn_normDist_T_656; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_658 = fmt0_recB_rawIn_fractIn[171] ? 9'h13c : _fmt0_recB_rawIn_normDist_T_657; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_659 = fmt0_recB_rawIn_fractIn[172] ? 9'h13b : _fmt0_recB_rawIn_normDist_T_658; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_660 = fmt0_recB_rawIn_fractIn[173] ? 9'h13a : _fmt0_recB_rawIn_normDist_T_659; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_661 = fmt0_recB_rawIn_fractIn[174] ? 9'h139 : _fmt0_recB_rawIn_normDist_T_660; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_662 = fmt0_recB_rawIn_fractIn[175] ? 9'h138 : _fmt0_recB_rawIn_normDist_T_661; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_663 = fmt0_recB_rawIn_fractIn[176] ? 9'h137 : _fmt0_recB_rawIn_normDist_T_662; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_664 = fmt0_recB_rawIn_fractIn[177] ? 9'h136 : _fmt0_recB_rawIn_normDist_T_663; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_665 = fmt0_recB_rawIn_fractIn[178] ? 9'h135 : _fmt0_recB_rawIn_normDist_T_664; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_666 = fmt0_recB_rawIn_fractIn[179] ? 9'h134 : _fmt0_recB_rawIn_normDist_T_665; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_667 = fmt0_recB_rawIn_fractIn[180] ? 9'h133 : _fmt0_recB_rawIn_normDist_T_666; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_668 = fmt0_recB_rawIn_fractIn[181] ? 9'h132 : _fmt0_recB_rawIn_normDist_T_667; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_669 = fmt0_recB_rawIn_fractIn[182] ? 9'h131 : _fmt0_recB_rawIn_normDist_T_668; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_670 = fmt0_recB_rawIn_fractIn[183] ? 9'h130 : _fmt0_recB_rawIn_normDist_T_669; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_671 = fmt0_recB_rawIn_fractIn[184] ? 9'h12f : _fmt0_recB_rawIn_normDist_T_670; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_672 = fmt0_recB_rawIn_fractIn[185] ? 9'h12e : _fmt0_recB_rawIn_normDist_T_671; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_673 = fmt0_recB_rawIn_fractIn[186] ? 9'h12d : _fmt0_recB_rawIn_normDist_T_672; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_674 = fmt0_recB_rawIn_fractIn[187] ? 9'h12c : _fmt0_recB_rawIn_normDist_T_673; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_675 = fmt0_recB_rawIn_fractIn[188] ? 9'h12b : _fmt0_recB_rawIn_normDist_T_674; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_676 = fmt0_recB_rawIn_fractIn[189] ? 9'h12a : _fmt0_recB_rawIn_normDist_T_675; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_677 = fmt0_recB_rawIn_fractIn[190] ? 9'h129 : _fmt0_recB_rawIn_normDist_T_676; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_678 = fmt0_recB_rawIn_fractIn[191] ? 9'h128 : _fmt0_recB_rawIn_normDist_T_677; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_679 = fmt0_recB_rawIn_fractIn[192] ? 9'h127 : _fmt0_recB_rawIn_normDist_T_678; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_680 = fmt0_recB_rawIn_fractIn[193] ? 9'h126 : _fmt0_recB_rawIn_normDist_T_679; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_681 = fmt0_recB_rawIn_fractIn[194] ? 9'h125 : _fmt0_recB_rawIn_normDist_T_680; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_682 = fmt0_recB_rawIn_fractIn[195] ? 9'h124 : _fmt0_recB_rawIn_normDist_T_681; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_683 = fmt0_recB_rawIn_fractIn[196] ? 9'h123 : _fmt0_recB_rawIn_normDist_T_682; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_684 = fmt0_recB_rawIn_fractIn[197] ? 9'h122 : _fmt0_recB_rawIn_normDist_T_683; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_685 = fmt0_recB_rawIn_fractIn[198] ? 9'h121 : _fmt0_recB_rawIn_normDist_T_684; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_686 = fmt0_recB_rawIn_fractIn[199] ? 9'h120 : _fmt0_recB_rawIn_normDist_T_685; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_687 = fmt0_recB_rawIn_fractIn[200] ? 9'h11f : _fmt0_recB_rawIn_normDist_T_686; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_688 = fmt0_recB_rawIn_fractIn[201] ? 9'h11e : _fmt0_recB_rawIn_normDist_T_687; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_689 = fmt0_recB_rawIn_fractIn[202] ? 9'h11d : _fmt0_recB_rawIn_normDist_T_688; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_690 = fmt0_recB_rawIn_fractIn[203] ? 9'h11c : _fmt0_recB_rawIn_normDist_T_689; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_691 = fmt0_recB_rawIn_fractIn[204] ? 9'h11b : _fmt0_recB_rawIn_normDist_T_690; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_692 = fmt0_recB_rawIn_fractIn[205] ? 9'h11a : _fmt0_recB_rawIn_normDist_T_691; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_693 = fmt0_recB_rawIn_fractIn[206] ? 9'h119 : _fmt0_recB_rawIn_normDist_T_692; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_694 = fmt0_recB_rawIn_fractIn[207] ? 9'h118 : _fmt0_recB_rawIn_normDist_T_693; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_695 = fmt0_recB_rawIn_fractIn[208] ? 9'h117 : _fmt0_recB_rawIn_normDist_T_694; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_696 = fmt0_recB_rawIn_fractIn[209] ? 9'h116 : _fmt0_recB_rawIn_normDist_T_695; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_697 = fmt0_recB_rawIn_fractIn[210] ? 9'h115 : _fmt0_recB_rawIn_normDist_T_696; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_698 = fmt0_recB_rawIn_fractIn[211] ? 9'h114 : _fmt0_recB_rawIn_normDist_T_697; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_699 = fmt0_recB_rawIn_fractIn[212] ? 9'h113 : _fmt0_recB_rawIn_normDist_T_698; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_700 = fmt0_recB_rawIn_fractIn[213] ? 9'h112 : _fmt0_recB_rawIn_normDist_T_699; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_701 = fmt0_recB_rawIn_fractIn[214] ? 9'h111 : _fmt0_recB_rawIn_normDist_T_700; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_702 = fmt0_recB_rawIn_fractIn[215] ? 9'h110 : _fmt0_recB_rawIn_normDist_T_701; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_703 = fmt0_recB_rawIn_fractIn[216] ? 9'h10f : _fmt0_recB_rawIn_normDist_T_702; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_704 = fmt0_recB_rawIn_fractIn[217] ? 9'h10e : _fmt0_recB_rawIn_normDist_T_703; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_705 = fmt0_recB_rawIn_fractIn[218] ? 9'h10d : _fmt0_recB_rawIn_normDist_T_704; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_706 = fmt0_recB_rawIn_fractIn[219] ? 9'h10c : _fmt0_recB_rawIn_normDist_T_705; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_707 = fmt0_recB_rawIn_fractIn[220] ? 9'h10b : _fmt0_recB_rawIn_normDist_T_706; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_708 = fmt0_recB_rawIn_fractIn[221] ? 9'h10a : _fmt0_recB_rawIn_normDist_T_707; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_709 = fmt0_recB_rawIn_fractIn[222] ? 9'h109 : _fmt0_recB_rawIn_normDist_T_708; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_710 = fmt0_recB_rawIn_fractIn[223] ? 9'h108 : _fmt0_recB_rawIn_normDist_T_709; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_711 = fmt0_recB_rawIn_fractIn[224] ? 9'h107 : _fmt0_recB_rawIn_normDist_T_710; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_712 = fmt0_recB_rawIn_fractIn[225] ? 9'h106 : _fmt0_recB_rawIn_normDist_T_711; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_713 = fmt0_recB_rawIn_fractIn[226] ? 9'h105 : _fmt0_recB_rawIn_normDist_T_712; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_714 = fmt0_recB_rawIn_fractIn[227] ? 9'h104 : _fmt0_recB_rawIn_normDist_T_713; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_715 = fmt0_recB_rawIn_fractIn[228] ? 9'h103 : _fmt0_recB_rawIn_normDist_T_714; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_716 = fmt0_recB_rawIn_fractIn[229] ? 9'h102 : _fmt0_recB_rawIn_normDist_T_715; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_717 = fmt0_recB_rawIn_fractIn[230] ? 9'h101 : _fmt0_recB_rawIn_normDist_T_716; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_718 = fmt0_recB_rawIn_fractIn[231] ? 9'h100 : _fmt0_recB_rawIn_normDist_T_717; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_719 = fmt0_recB_rawIn_fractIn[232] ? 9'hff : _fmt0_recB_rawIn_normDist_T_718; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_720 = fmt0_recB_rawIn_fractIn[233] ? 9'hfe : _fmt0_recB_rawIn_normDist_T_719; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_721 = fmt0_recB_rawIn_fractIn[234] ? 9'hfd : _fmt0_recB_rawIn_normDist_T_720; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_722 = fmt0_recB_rawIn_fractIn[235] ? 9'hfc : _fmt0_recB_rawIn_normDist_T_721; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_723 = fmt0_recB_rawIn_fractIn[236] ? 9'hfb : _fmt0_recB_rawIn_normDist_T_722; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_724 = fmt0_recB_rawIn_fractIn[237] ? 9'hfa : _fmt0_recB_rawIn_normDist_T_723; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_725 = fmt0_recB_rawIn_fractIn[238] ? 9'hf9 : _fmt0_recB_rawIn_normDist_T_724; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_726 = fmt0_recB_rawIn_fractIn[239] ? 9'hf8 : _fmt0_recB_rawIn_normDist_T_725; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_727 = fmt0_recB_rawIn_fractIn[240] ? 9'hf7 : _fmt0_recB_rawIn_normDist_T_726; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_728 = fmt0_recB_rawIn_fractIn[241] ? 9'hf6 : _fmt0_recB_rawIn_normDist_T_727; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_729 = fmt0_recB_rawIn_fractIn[242] ? 9'hf5 : _fmt0_recB_rawIn_normDist_T_728; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_730 = fmt0_recB_rawIn_fractIn[243] ? 9'hf4 : _fmt0_recB_rawIn_normDist_T_729; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_731 = fmt0_recB_rawIn_fractIn[244] ? 9'hf3 : _fmt0_recB_rawIn_normDist_T_730; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_732 = fmt0_recB_rawIn_fractIn[245] ? 9'hf2 : _fmt0_recB_rawIn_normDist_T_731; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_733 = fmt0_recB_rawIn_fractIn[246] ? 9'hf1 : _fmt0_recB_rawIn_normDist_T_732; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_734 = fmt0_recB_rawIn_fractIn[247] ? 9'hf0 : _fmt0_recB_rawIn_normDist_T_733; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_735 = fmt0_recB_rawIn_fractIn[248] ? 9'hef : _fmt0_recB_rawIn_normDist_T_734; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_736 = fmt0_recB_rawIn_fractIn[249] ? 9'hee : _fmt0_recB_rawIn_normDist_T_735; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_737 = fmt0_recB_rawIn_fractIn[250] ? 9'hed : _fmt0_recB_rawIn_normDist_T_736; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_738 = fmt0_recB_rawIn_fractIn[251] ? 9'hec : _fmt0_recB_rawIn_normDist_T_737; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_739 = fmt0_recB_rawIn_fractIn[252] ? 9'heb : _fmt0_recB_rawIn_normDist_T_738; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_740 = fmt0_recB_rawIn_fractIn[253] ? 9'hea : _fmt0_recB_rawIn_normDist_T_739; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_741 = fmt0_recB_rawIn_fractIn[254] ? 9'he9 : _fmt0_recB_rawIn_normDist_T_740; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_742 = fmt0_recB_rawIn_fractIn[255] ? 9'he8 : _fmt0_recB_rawIn_normDist_T_741; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_743 = fmt0_recB_rawIn_fractIn[256] ? 9'he7 : _fmt0_recB_rawIn_normDist_T_742; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_744 = fmt0_recB_rawIn_fractIn[257] ? 9'he6 : _fmt0_recB_rawIn_normDist_T_743; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_745 = fmt0_recB_rawIn_fractIn[258] ? 9'he5 : _fmt0_recB_rawIn_normDist_T_744; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_746 = fmt0_recB_rawIn_fractIn[259] ? 9'he4 : _fmt0_recB_rawIn_normDist_T_745; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_747 = fmt0_recB_rawIn_fractIn[260] ? 9'he3 : _fmt0_recB_rawIn_normDist_T_746; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_748 = fmt0_recB_rawIn_fractIn[261] ? 9'he2 : _fmt0_recB_rawIn_normDist_T_747; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_749 = fmt0_recB_rawIn_fractIn[262] ? 9'he1 : _fmt0_recB_rawIn_normDist_T_748; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_750 = fmt0_recB_rawIn_fractIn[263] ? 9'he0 : _fmt0_recB_rawIn_normDist_T_749; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_751 = fmt0_recB_rawIn_fractIn[264] ? 9'hdf : _fmt0_recB_rawIn_normDist_T_750; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_752 = fmt0_recB_rawIn_fractIn[265] ? 9'hde : _fmt0_recB_rawIn_normDist_T_751; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_753 = fmt0_recB_rawIn_fractIn[266] ? 9'hdd : _fmt0_recB_rawIn_normDist_T_752; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_754 = fmt0_recB_rawIn_fractIn[267] ? 9'hdc : _fmt0_recB_rawIn_normDist_T_753; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_755 = fmt0_recB_rawIn_fractIn[268] ? 9'hdb : _fmt0_recB_rawIn_normDist_T_754; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_756 = fmt0_recB_rawIn_fractIn[269] ? 9'hda : _fmt0_recB_rawIn_normDist_T_755; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_757 = fmt0_recB_rawIn_fractIn[270] ? 9'hd9 : _fmt0_recB_rawIn_normDist_T_756; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_758 = fmt0_recB_rawIn_fractIn[271] ? 9'hd8 : _fmt0_recB_rawIn_normDist_T_757; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_759 = fmt0_recB_rawIn_fractIn[272] ? 9'hd7 : _fmt0_recB_rawIn_normDist_T_758; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_760 = fmt0_recB_rawIn_fractIn[273] ? 9'hd6 : _fmt0_recB_rawIn_normDist_T_759; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_761 = fmt0_recB_rawIn_fractIn[274] ? 9'hd5 : _fmt0_recB_rawIn_normDist_T_760; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_762 = fmt0_recB_rawIn_fractIn[275] ? 9'hd4 : _fmt0_recB_rawIn_normDist_T_761; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_763 = fmt0_recB_rawIn_fractIn[276] ? 9'hd3 : _fmt0_recB_rawIn_normDist_T_762; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_764 = fmt0_recB_rawIn_fractIn[277] ? 9'hd2 : _fmt0_recB_rawIn_normDist_T_763; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_765 = fmt0_recB_rawIn_fractIn[278] ? 9'hd1 : _fmt0_recB_rawIn_normDist_T_764; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_766 = fmt0_recB_rawIn_fractIn[279] ? 9'hd0 : _fmt0_recB_rawIn_normDist_T_765; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_767 = fmt0_recB_rawIn_fractIn[280] ? 9'hcf : _fmt0_recB_rawIn_normDist_T_766; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_768 = fmt0_recB_rawIn_fractIn[281] ? 9'hce : _fmt0_recB_rawIn_normDist_T_767; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_769 = fmt0_recB_rawIn_fractIn[282] ? 9'hcd : _fmt0_recB_rawIn_normDist_T_768; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_770 = fmt0_recB_rawIn_fractIn[283] ? 9'hcc : _fmt0_recB_rawIn_normDist_T_769; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_771 = fmt0_recB_rawIn_fractIn[284] ? 9'hcb : _fmt0_recB_rawIn_normDist_T_770; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_772 = fmt0_recB_rawIn_fractIn[285] ? 9'hca : _fmt0_recB_rawIn_normDist_T_771; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_773 = fmt0_recB_rawIn_fractIn[286] ? 9'hc9 : _fmt0_recB_rawIn_normDist_T_772; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_774 = fmt0_recB_rawIn_fractIn[287] ? 9'hc8 : _fmt0_recB_rawIn_normDist_T_773; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_775 = fmt0_recB_rawIn_fractIn[288] ? 9'hc7 : _fmt0_recB_rawIn_normDist_T_774; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_776 = fmt0_recB_rawIn_fractIn[289] ? 9'hc6 : _fmt0_recB_rawIn_normDist_T_775; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_777 = fmt0_recB_rawIn_fractIn[290] ? 9'hc5 : _fmt0_recB_rawIn_normDist_T_776; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_778 = fmt0_recB_rawIn_fractIn[291] ? 9'hc4 : _fmt0_recB_rawIn_normDist_T_777; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_779 = fmt0_recB_rawIn_fractIn[292] ? 9'hc3 : _fmt0_recB_rawIn_normDist_T_778; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_780 = fmt0_recB_rawIn_fractIn[293] ? 9'hc2 : _fmt0_recB_rawIn_normDist_T_779; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_781 = fmt0_recB_rawIn_fractIn[294] ? 9'hc1 : _fmt0_recB_rawIn_normDist_T_780; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_782 = fmt0_recB_rawIn_fractIn[295] ? 9'hc0 : _fmt0_recB_rawIn_normDist_T_781; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_783 = fmt0_recB_rawIn_fractIn[296] ? 9'hbf : _fmt0_recB_rawIn_normDist_T_782; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_784 = fmt0_recB_rawIn_fractIn[297] ? 9'hbe : _fmt0_recB_rawIn_normDist_T_783; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_785 = fmt0_recB_rawIn_fractIn[298] ? 9'hbd : _fmt0_recB_rawIn_normDist_T_784; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_786 = fmt0_recB_rawIn_fractIn[299] ? 9'hbc : _fmt0_recB_rawIn_normDist_T_785; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_787 = fmt0_recB_rawIn_fractIn[300] ? 9'hbb : _fmt0_recB_rawIn_normDist_T_786; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_788 = fmt0_recB_rawIn_fractIn[301] ? 9'hba : _fmt0_recB_rawIn_normDist_T_787; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_789 = fmt0_recB_rawIn_fractIn[302] ? 9'hb9 : _fmt0_recB_rawIn_normDist_T_788; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_790 = fmt0_recB_rawIn_fractIn[303] ? 9'hb8 : _fmt0_recB_rawIn_normDist_T_789; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_791 = fmt0_recB_rawIn_fractIn[304] ? 9'hb7 : _fmt0_recB_rawIn_normDist_T_790; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_792 = fmt0_recB_rawIn_fractIn[305] ? 9'hb6 : _fmt0_recB_rawIn_normDist_T_791; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_793 = fmt0_recB_rawIn_fractIn[306] ? 9'hb5 : _fmt0_recB_rawIn_normDist_T_792; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_794 = fmt0_recB_rawIn_fractIn[307] ? 9'hb4 : _fmt0_recB_rawIn_normDist_T_793; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_795 = fmt0_recB_rawIn_fractIn[308] ? 9'hb3 : _fmt0_recB_rawIn_normDist_T_794; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_796 = fmt0_recB_rawIn_fractIn[309] ? 9'hb2 : _fmt0_recB_rawIn_normDist_T_795; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_797 = fmt0_recB_rawIn_fractIn[310] ? 9'hb1 : _fmt0_recB_rawIn_normDist_T_796; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_798 = fmt0_recB_rawIn_fractIn[311] ? 9'hb0 : _fmt0_recB_rawIn_normDist_T_797; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_799 = fmt0_recB_rawIn_fractIn[312] ? 9'haf : _fmt0_recB_rawIn_normDist_T_798; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_800 = fmt0_recB_rawIn_fractIn[313] ? 9'hae : _fmt0_recB_rawIn_normDist_T_799; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_801 = fmt0_recB_rawIn_fractIn[314] ? 9'had : _fmt0_recB_rawIn_normDist_T_800; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_802 = fmt0_recB_rawIn_fractIn[315] ? 9'hac : _fmt0_recB_rawIn_normDist_T_801; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_803 = fmt0_recB_rawIn_fractIn[316] ? 9'hab : _fmt0_recB_rawIn_normDist_T_802; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_804 = fmt0_recB_rawIn_fractIn[317] ? 9'haa : _fmt0_recB_rawIn_normDist_T_803; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_805 = fmt0_recB_rawIn_fractIn[318] ? 9'ha9 : _fmt0_recB_rawIn_normDist_T_804; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_806 = fmt0_recB_rawIn_fractIn[319] ? 9'ha8 : _fmt0_recB_rawIn_normDist_T_805; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_807 = fmt0_recB_rawIn_fractIn[320] ? 9'ha7 : _fmt0_recB_rawIn_normDist_T_806; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_808 = fmt0_recB_rawIn_fractIn[321] ? 9'ha6 : _fmt0_recB_rawIn_normDist_T_807; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_809 = fmt0_recB_rawIn_fractIn[322] ? 9'ha5 : _fmt0_recB_rawIn_normDist_T_808; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_810 = fmt0_recB_rawIn_fractIn[323] ? 9'ha4 : _fmt0_recB_rawIn_normDist_T_809; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_811 = fmt0_recB_rawIn_fractIn[324] ? 9'ha3 : _fmt0_recB_rawIn_normDist_T_810; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_812 = fmt0_recB_rawIn_fractIn[325] ? 9'ha2 : _fmt0_recB_rawIn_normDist_T_811; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_813 = fmt0_recB_rawIn_fractIn[326] ? 9'ha1 : _fmt0_recB_rawIn_normDist_T_812; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_814 = fmt0_recB_rawIn_fractIn[327] ? 9'ha0 : _fmt0_recB_rawIn_normDist_T_813; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_815 = fmt0_recB_rawIn_fractIn[328] ? 9'h9f : _fmt0_recB_rawIn_normDist_T_814; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_816 = fmt0_recB_rawIn_fractIn[329] ? 9'h9e : _fmt0_recB_rawIn_normDist_T_815; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_817 = fmt0_recB_rawIn_fractIn[330] ? 9'h9d : _fmt0_recB_rawIn_normDist_T_816; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_818 = fmt0_recB_rawIn_fractIn[331] ? 9'h9c : _fmt0_recB_rawIn_normDist_T_817; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_819 = fmt0_recB_rawIn_fractIn[332] ? 9'h9b : _fmt0_recB_rawIn_normDist_T_818; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_820 = fmt0_recB_rawIn_fractIn[333] ? 9'h9a : _fmt0_recB_rawIn_normDist_T_819; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_821 = fmt0_recB_rawIn_fractIn[334] ? 9'h99 : _fmt0_recB_rawIn_normDist_T_820; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_822 = fmt0_recB_rawIn_fractIn[335] ? 9'h98 : _fmt0_recB_rawIn_normDist_T_821; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_823 = fmt0_recB_rawIn_fractIn[336] ? 9'h97 : _fmt0_recB_rawIn_normDist_T_822; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_824 = fmt0_recB_rawIn_fractIn[337] ? 9'h96 : _fmt0_recB_rawIn_normDist_T_823; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_825 = fmt0_recB_rawIn_fractIn[338] ? 9'h95 : _fmt0_recB_rawIn_normDist_T_824; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_826 = fmt0_recB_rawIn_fractIn[339] ? 9'h94 : _fmt0_recB_rawIn_normDist_T_825; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_827 = fmt0_recB_rawIn_fractIn[340] ? 9'h93 : _fmt0_recB_rawIn_normDist_T_826; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_828 = fmt0_recB_rawIn_fractIn[341] ? 9'h92 : _fmt0_recB_rawIn_normDist_T_827; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_829 = fmt0_recB_rawIn_fractIn[342] ? 9'h91 : _fmt0_recB_rawIn_normDist_T_828; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_830 = fmt0_recB_rawIn_fractIn[343] ? 9'h90 : _fmt0_recB_rawIn_normDist_T_829; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_831 = fmt0_recB_rawIn_fractIn[344] ? 9'h8f : _fmt0_recB_rawIn_normDist_T_830; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_832 = fmt0_recB_rawIn_fractIn[345] ? 9'h8e : _fmt0_recB_rawIn_normDist_T_831; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_833 = fmt0_recB_rawIn_fractIn[346] ? 9'h8d : _fmt0_recB_rawIn_normDist_T_832; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_834 = fmt0_recB_rawIn_fractIn[347] ? 9'h8c : _fmt0_recB_rawIn_normDist_T_833; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_835 = fmt0_recB_rawIn_fractIn[348] ? 9'h8b : _fmt0_recB_rawIn_normDist_T_834; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_836 = fmt0_recB_rawIn_fractIn[349] ? 9'h8a : _fmt0_recB_rawIn_normDist_T_835; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_837 = fmt0_recB_rawIn_fractIn[350] ? 9'h89 : _fmt0_recB_rawIn_normDist_T_836; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_838 = fmt0_recB_rawIn_fractIn[351] ? 9'h88 : _fmt0_recB_rawIn_normDist_T_837; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_839 = fmt0_recB_rawIn_fractIn[352] ? 9'h87 : _fmt0_recB_rawIn_normDist_T_838; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_840 = fmt0_recB_rawIn_fractIn[353] ? 9'h86 : _fmt0_recB_rawIn_normDist_T_839; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_841 = fmt0_recB_rawIn_fractIn[354] ? 9'h85 : _fmt0_recB_rawIn_normDist_T_840; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_842 = fmt0_recB_rawIn_fractIn[355] ? 9'h84 : _fmt0_recB_rawIn_normDist_T_841; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_843 = fmt0_recB_rawIn_fractIn[356] ? 9'h83 : _fmt0_recB_rawIn_normDist_T_842; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_844 = fmt0_recB_rawIn_fractIn[357] ? 9'h82 : _fmt0_recB_rawIn_normDist_T_843; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_845 = fmt0_recB_rawIn_fractIn[358] ? 9'h81 : _fmt0_recB_rawIn_normDist_T_844; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_846 = fmt0_recB_rawIn_fractIn[359] ? 9'h80 : _fmt0_recB_rawIn_normDist_T_845; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_847 = fmt0_recB_rawIn_fractIn[360] ? 9'h7f : _fmt0_recB_rawIn_normDist_T_846; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_848 = fmt0_recB_rawIn_fractIn[361] ? 9'h7e : _fmt0_recB_rawIn_normDist_T_847; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_849 = fmt0_recB_rawIn_fractIn[362] ? 9'h7d : _fmt0_recB_rawIn_normDist_T_848; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_850 = fmt0_recB_rawIn_fractIn[363] ? 9'h7c : _fmt0_recB_rawIn_normDist_T_849; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_851 = fmt0_recB_rawIn_fractIn[364] ? 9'h7b : _fmt0_recB_rawIn_normDist_T_850; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_852 = fmt0_recB_rawIn_fractIn[365] ? 9'h7a : _fmt0_recB_rawIn_normDist_T_851; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_853 = fmt0_recB_rawIn_fractIn[366] ? 9'h79 : _fmt0_recB_rawIn_normDist_T_852; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_854 = fmt0_recB_rawIn_fractIn[367] ? 9'h78 : _fmt0_recB_rawIn_normDist_T_853; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_855 = fmt0_recB_rawIn_fractIn[368] ? 9'h77 : _fmt0_recB_rawIn_normDist_T_854; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_856 = fmt0_recB_rawIn_fractIn[369] ? 9'h76 : _fmt0_recB_rawIn_normDist_T_855; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_857 = fmt0_recB_rawIn_fractIn[370] ? 9'h75 : _fmt0_recB_rawIn_normDist_T_856; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_858 = fmt0_recB_rawIn_fractIn[371] ? 9'h74 : _fmt0_recB_rawIn_normDist_T_857; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_859 = fmt0_recB_rawIn_fractIn[372] ? 9'h73 : _fmt0_recB_rawIn_normDist_T_858; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_860 = fmt0_recB_rawIn_fractIn[373] ? 9'h72 : _fmt0_recB_rawIn_normDist_T_859; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_861 = fmt0_recB_rawIn_fractIn[374] ? 9'h71 : _fmt0_recB_rawIn_normDist_T_860; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_862 = fmt0_recB_rawIn_fractIn[375] ? 9'h70 : _fmt0_recB_rawIn_normDist_T_861; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_863 = fmt0_recB_rawIn_fractIn[376] ? 9'h6f : _fmt0_recB_rawIn_normDist_T_862; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_864 = fmt0_recB_rawIn_fractIn[377] ? 9'h6e : _fmt0_recB_rawIn_normDist_T_863; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_865 = fmt0_recB_rawIn_fractIn[378] ? 9'h6d : _fmt0_recB_rawIn_normDist_T_864; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_866 = fmt0_recB_rawIn_fractIn[379] ? 9'h6c : _fmt0_recB_rawIn_normDist_T_865; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_867 = fmt0_recB_rawIn_fractIn[380] ? 9'h6b : _fmt0_recB_rawIn_normDist_T_866; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_868 = fmt0_recB_rawIn_fractIn[381] ? 9'h6a : _fmt0_recB_rawIn_normDist_T_867; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_869 = fmt0_recB_rawIn_fractIn[382] ? 9'h69 : _fmt0_recB_rawIn_normDist_T_868; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_870 = fmt0_recB_rawIn_fractIn[383] ? 9'h68 : _fmt0_recB_rawIn_normDist_T_869; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_871 = fmt0_recB_rawIn_fractIn[384] ? 9'h67 : _fmt0_recB_rawIn_normDist_T_870; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_872 = fmt0_recB_rawIn_fractIn[385] ? 9'h66 : _fmt0_recB_rawIn_normDist_T_871; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_873 = fmt0_recB_rawIn_fractIn[386] ? 9'h65 : _fmt0_recB_rawIn_normDist_T_872; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_874 = fmt0_recB_rawIn_fractIn[387] ? 9'h64 : _fmt0_recB_rawIn_normDist_T_873; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_875 = fmt0_recB_rawIn_fractIn[388] ? 9'h63 : _fmt0_recB_rawIn_normDist_T_874; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_876 = fmt0_recB_rawIn_fractIn[389] ? 9'h62 : _fmt0_recB_rawIn_normDist_T_875; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_877 = fmt0_recB_rawIn_fractIn[390] ? 9'h61 : _fmt0_recB_rawIn_normDist_T_876; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_878 = fmt0_recB_rawIn_fractIn[391] ? 9'h60 : _fmt0_recB_rawIn_normDist_T_877; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_879 = fmt0_recB_rawIn_fractIn[392] ? 9'h5f : _fmt0_recB_rawIn_normDist_T_878; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_880 = fmt0_recB_rawIn_fractIn[393] ? 9'h5e : _fmt0_recB_rawIn_normDist_T_879; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_881 = fmt0_recB_rawIn_fractIn[394] ? 9'h5d : _fmt0_recB_rawIn_normDist_T_880; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_882 = fmt0_recB_rawIn_fractIn[395] ? 9'h5c : _fmt0_recB_rawIn_normDist_T_881; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_883 = fmt0_recB_rawIn_fractIn[396] ? 9'h5b : _fmt0_recB_rawIn_normDist_T_882; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_884 = fmt0_recB_rawIn_fractIn[397] ? 9'h5a : _fmt0_recB_rawIn_normDist_T_883; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_885 = fmt0_recB_rawIn_fractIn[398] ? 9'h59 : _fmt0_recB_rawIn_normDist_T_884; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_886 = fmt0_recB_rawIn_fractIn[399] ? 9'h58 : _fmt0_recB_rawIn_normDist_T_885; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_887 = fmt0_recB_rawIn_fractIn[400] ? 9'h57 : _fmt0_recB_rawIn_normDist_T_886; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_888 = fmt0_recB_rawIn_fractIn[401] ? 9'h56 : _fmt0_recB_rawIn_normDist_T_887; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_889 = fmt0_recB_rawIn_fractIn[402] ? 9'h55 : _fmt0_recB_rawIn_normDist_T_888; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_890 = fmt0_recB_rawIn_fractIn[403] ? 9'h54 : _fmt0_recB_rawIn_normDist_T_889; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_891 = fmt0_recB_rawIn_fractIn[404] ? 9'h53 : _fmt0_recB_rawIn_normDist_T_890; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_892 = fmt0_recB_rawIn_fractIn[405] ? 9'h52 : _fmt0_recB_rawIn_normDist_T_891; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_893 = fmt0_recB_rawIn_fractIn[406] ? 9'h51 : _fmt0_recB_rawIn_normDist_T_892; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_894 = fmt0_recB_rawIn_fractIn[407] ? 9'h50 : _fmt0_recB_rawIn_normDist_T_893; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_895 = fmt0_recB_rawIn_fractIn[408] ? 9'h4f : _fmt0_recB_rawIn_normDist_T_894; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_896 = fmt0_recB_rawIn_fractIn[409] ? 9'h4e : _fmt0_recB_rawIn_normDist_T_895; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_897 = fmt0_recB_rawIn_fractIn[410] ? 9'h4d : _fmt0_recB_rawIn_normDist_T_896; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_898 = fmt0_recB_rawIn_fractIn[411] ? 9'h4c : _fmt0_recB_rawIn_normDist_T_897; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_899 = fmt0_recB_rawIn_fractIn[412] ? 9'h4b : _fmt0_recB_rawIn_normDist_T_898; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_900 = fmt0_recB_rawIn_fractIn[413] ? 9'h4a : _fmt0_recB_rawIn_normDist_T_899; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_901 = fmt0_recB_rawIn_fractIn[414] ? 9'h49 : _fmt0_recB_rawIn_normDist_T_900; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_902 = fmt0_recB_rawIn_fractIn[415] ? 9'h48 : _fmt0_recB_rawIn_normDist_T_901; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_903 = fmt0_recB_rawIn_fractIn[416] ? 9'h47 : _fmt0_recB_rawIn_normDist_T_902; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_904 = fmt0_recB_rawIn_fractIn[417] ? 9'h46 : _fmt0_recB_rawIn_normDist_T_903; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_905 = fmt0_recB_rawIn_fractIn[418] ? 9'h45 : _fmt0_recB_rawIn_normDist_T_904; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_906 = fmt0_recB_rawIn_fractIn[419] ? 9'h44 : _fmt0_recB_rawIn_normDist_T_905; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_907 = fmt0_recB_rawIn_fractIn[420] ? 9'h43 : _fmt0_recB_rawIn_normDist_T_906; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_908 = fmt0_recB_rawIn_fractIn[421] ? 9'h42 : _fmt0_recB_rawIn_normDist_T_907; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_909 = fmt0_recB_rawIn_fractIn[422] ? 9'h41 : _fmt0_recB_rawIn_normDist_T_908; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_910 = fmt0_recB_rawIn_fractIn[423] ? 9'h40 : _fmt0_recB_rawIn_normDist_T_909; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_911 = fmt0_recB_rawIn_fractIn[424] ? 9'h3f : _fmt0_recB_rawIn_normDist_T_910; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_912 = fmt0_recB_rawIn_fractIn[425] ? 9'h3e : _fmt0_recB_rawIn_normDist_T_911; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_913 = fmt0_recB_rawIn_fractIn[426] ? 9'h3d : _fmt0_recB_rawIn_normDist_T_912; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_914 = fmt0_recB_rawIn_fractIn[427] ? 9'h3c : _fmt0_recB_rawIn_normDist_T_913; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_915 = fmt0_recB_rawIn_fractIn[428] ? 9'h3b : _fmt0_recB_rawIn_normDist_T_914; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_916 = fmt0_recB_rawIn_fractIn[429] ? 9'h3a : _fmt0_recB_rawIn_normDist_T_915; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_917 = fmt0_recB_rawIn_fractIn[430] ? 9'h39 : _fmt0_recB_rawIn_normDist_T_916; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_918 = fmt0_recB_rawIn_fractIn[431] ? 9'h38 : _fmt0_recB_rawIn_normDist_T_917; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_919 = fmt0_recB_rawIn_fractIn[432] ? 9'h37 : _fmt0_recB_rawIn_normDist_T_918; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_920 = fmt0_recB_rawIn_fractIn[433] ? 9'h36 : _fmt0_recB_rawIn_normDist_T_919; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_921 = fmt0_recB_rawIn_fractIn[434] ? 9'h35 : _fmt0_recB_rawIn_normDist_T_920; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_922 = fmt0_recB_rawIn_fractIn[435] ? 9'h34 : _fmt0_recB_rawIn_normDist_T_921; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_923 = fmt0_recB_rawIn_fractIn[436] ? 9'h33 : _fmt0_recB_rawIn_normDist_T_922; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_924 = fmt0_recB_rawIn_fractIn[437] ? 9'h32 : _fmt0_recB_rawIn_normDist_T_923; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_925 = fmt0_recB_rawIn_fractIn[438] ? 9'h31 : _fmt0_recB_rawIn_normDist_T_924; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_926 = fmt0_recB_rawIn_fractIn[439] ? 9'h30 : _fmt0_recB_rawIn_normDist_T_925; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_927 = fmt0_recB_rawIn_fractIn[440] ? 9'h2f : _fmt0_recB_rawIn_normDist_T_926; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_928 = fmt0_recB_rawIn_fractIn[441] ? 9'h2e : _fmt0_recB_rawIn_normDist_T_927; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_929 = fmt0_recB_rawIn_fractIn[442] ? 9'h2d : _fmt0_recB_rawIn_normDist_T_928; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_930 = fmt0_recB_rawIn_fractIn[443] ? 9'h2c : _fmt0_recB_rawIn_normDist_T_929; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_931 = fmt0_recB_rawIn_fractIn[444] ? 9'h2b : _fmt0_recB_rawIn_normDist_T_930; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_932 = fmt0_recB_rawIn_fractIn[445] ? 9'h2a : _fmt0_recB_rawIn_normDist_T_931; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_933 = fmt0_recB_rawIn_fractIn[446] ? 9'h29 : _fmt0_recB_rawIn_normDist_T_932; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_934 = fmt0_recB_rawIn_fractIn[447] ? 9'h28 : _fmt0_recB_rawIn_normDist_T_933; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_935 = fmt0_recB_rawIn_fractIn[448] ? 9'h27 : _fmt0_recB_rawIn_normDist_T_934; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_936 = fmt0_recB_rawIn_fractIn[449] ? 9'h26 : _fmt0_recB_rawIn_normDist_T_935; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_937 = fmt0_recB_rawIn_fractIn[450] ? 9'h25 : _fmt0_recB_rawIn_normDist_T_936; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_938 = fmt0_recB_rawIn_fractIn[451] ? 9'h24 : _fmt0_recB_rawIn_normDist_T_937; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_939 = fmt0_recB_rawIn_fractIn[452] ? 9'h23 : _fmt0_recB_rawIn_normDist_T_938; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_940 = fmt0_recB_rawIn_fractIn[453] ? 9'h22 : _fmt0_recB_rawIn_normDist_T_939; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_941 = fmt0_recB_rawIn_fractIn[454] ? 9'h21 : _fmt0_recB_rawIn_normDist_T_940; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_942 = fmt0_recB_rawIn_fractIn[455] ? 9'h20 : _fmt0_recB_rawIn_normDist_T_941; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_943 = fmt0_recB_rawIn_fractIn[456] ? 9'h1f : _fmt0_recB_rawIn_normDist_T_942; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_944 = fmt0_recB_rawIn_fractIn[457] ? 9'h1e : _fmt0_recB_rawIn_normDist_T_943; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_945 = fmt0_recB_rawIn_fractIn[458] ? 9'h1d : _fmt0_recB_rawIn_normDist_T_944; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_946 = fmt0_recB_rawIn_fractIn[459] ? 9'h1c : _fmt0_recB_rawIn_normDist_T_945; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_947 = fmt0_recB_rawIn_fractIn[460] ? 9'h1b : _fmt0_recB_rawIn_normDist_T_946; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_948 = fmt0_recB_rawIn_fractIn[461] ? 9'h1a : _fmt0_recB_rawIn_normDist_T_947; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_949 = fmt0_recB_rawIn_fractIn[462] ? 9'h19 : _fmt0_recB_rawIn_normDist_T_948; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_950 = fmt0_recB_rawIn_fractIn[463] ? 9'h18 : _fmt0_recB_rawIn_normDist_T_949; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_951 = fmt0_recB_rawIn_fractIn[464] ? 9'h17 : _fmt0_recB_rawIn_normDist_T_950; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_952 = fmt0_recB_rawIn_fractIn[465] ? 9'h16 : _fmt0_recB_rawIn_normDist_T_951; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_953 = fmt0_recB_rawIn_fractIn[466] ? 9'h15 : _fmt0_recB_rawIn_normDist_T_952; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_954 = fmt0_recB_rawIn_fractIn[467] ? 9'h14 : _fmt0_recB_rawIn_normDist_T_953; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_955 = fmt0_recB_rawIn_fractIn[468] ? 9'h13 : _fmt0_recB_rawIn_normDist_T_954; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_956 = fmt0_recB_rawIn_fractIn[469] ? 9'h12 : _fmt0_recB_rawIn_normDist_T_955; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_957 = fmt0_recB_rawIn_fractIn[470] ? 9'h11 : _fmt0_recB_rawIn_normDist_T_956; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_958 = fmt0_recB_rawIn_fractIn[471] ? 9'h10 : _fmt0_recB_rawIn_normDist_T_957; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_959 = fmt0_recB_rawIn_fractIn[472] ? 9'hf : _fmt0_recB_rawIn_normDist_T_958; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_960 = fmt0_recB_rawIn_fractIn[473] ? 9'he : _fmt0_recB_rawIn_normDist_T_959; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_961 = fmt0_recB_rawIn_fractIn[474] ? 9'hd : _fmt0_recB_rawIn_normDist_T_960; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_962 = fmt0_recB_rawIn_fractIn[475] ? 9'hc : _fmt0_recB_rawIn_normDist_T_961; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_963 = fmt0_recB_rawIn_fractIn[476] ? 9'hb : _fmt0_recB_rawIn_normDist_T_962; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_964 = fmt0_recB_rawIn_fractIn[477] ? 9'ha : _fmt0_recB_rawIn_normDist_T_963; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_965 = fmt0_recB_rawIn_fractIn[478] ? 9'h9 : _fmt0_recB_rawIn_normDist_T_964; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_966 = fmt0_recB_rawIn_fractIn[479] ? 9'h8 : _fmt0_recB_rawIn_normDist_T_965; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_967 = fmt0_recB_rawIn_fractIn[480] ? 9'h7 : _fmt0_recB_rawIn_normDist_T_966; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_968 = fmt0_recB_rawIn_fractIn[481] ? 9'h6 : _fmt0_recB_rawIn_normDist_T_967; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_969 = fmt0_recB_rawIn_fractIn[482] ? 9'h5 : _fmt0_recB_rawIn_normDist_T_968; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_970 = fmt0_recB_rawIn_fractIn[483] ? 9'h4 : _fmt0_recB_rawIn_normDist_T_969; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_971 = fmt0_recB_rawIn_fractIn[484] ? 9'h3 : _fmt0_recB_rawIn_normDist_T_970; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_972 = fmt0_recB_rawIn_fractIn[485] ? 9'h2 : _fmt0_recB_rawIn_normDist_T_971; // @[Mux.scala 47:70]
  wire [8:0] _fmt0_recB_rawIn_normDist_T_973 = fmt0_recB_rawIn_fractIn[486] ? 9'h1 : _fmt0_recB_rawIn_normDist_T_972; // @[Mux.scala 47:70]
  wire [8:0] fmt0_recB_rawIn_normDist = fmt0_recB_rawIn_fractIn[487] ? 9'h0 : _fmt0_recB_rawIn_normDist_T_973; // @[Mux.scala 47:70]
  wire [998:0] _GEN_6 = {{511'd0}, fmt0_recB_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [998:0] _fmt0_recB_rawIn_subnormFract_T = _GEN_6 << fmt0_recB_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [487:0] fmt0_recB_rawIn_subnormFract = {_fmt0_recB_rawIn_subnormFract_T[486:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [23:0] _GEN_13 = {{15'd0}, fmt0_recB_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [23:0] _fmt0_recB_rawIn_adjustedExp_T = _GEN_13 ^ 24'hffffff; // @[rawFloatFromFN.scala 55:18]
  wire [23:0] _fmt0_recB_rawIn_adjustedExp_T_1 = fmt0_recB_rawIn_isZeroExpIn ? _fmt0_recB_rawIn_adjustedExp_T : {{1
    'd0}, fmt0_recB_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _fmt0_recB_rawIn_adjustedExp_T_2 = fmt0_recB_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [22:0] _GEN_14 = {{21'd0}, _fmt0_recB_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [22:0] _fmt0_recB_rawIn_adjustedExp_T_3 = 23'h400000 | _GEN_14; // @[rawFloatFromFN.scala 58:9]
  wire [23:0] _GEN_15 = {{1'd0}, _fmt0_recB_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [23:0] fmt0_recB_rawIn_adjustedExp = _fmt0_recB_rawIn_adjustedExp_T_1 + _GEN_15; // @[rawFloatFromFN.scala 57:9]
  wire  fmt0_recB_rawIn_isZero = fmt0_recB_rawIn_isZeroExpIn & fmt0_recB_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  fmt0_recB_rawIn_isSpecial = fmt0_recB_rawIn_adjustedExp[23:22] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  fmt0_recB_rawIn__isNaN = fmt0_recB_rawIn_isSpecial & ~fmt0_recB_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [24:0] fmt0_recB_rawIn__sExp = {1'b0,$signed(fmt0_recB_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _fmt0_recB_rawIn_out_sig_T = ~fmt0_recB_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [487:0] _fmt0_recB_rawIn_out_sig_T_2 = fmt0_recB_rawIn_isZeroExpIn ? fmt0_recB_rawIn_subnormFract :
    fmt0_recB_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [489:0] fmt0_recB_rawIn__sig = {1'h0,_fmt0_recB_rawIn_out_sig_T,_fmt0_recB_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _fmt0_recB_T_2 = fmt0_recB_rawIn_isZero ? 3'h0 : fmt0_recB_rawIn__sExp[23:21]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_16 = {{2'd0}, fmt0_recB_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _fmt0_recB_T_4 = _fmt0_recB_T_2 | _GEN_16; // @[recFNFromFN.scala 48:76]
  wire [24:0] _fmt0_recB_T_7 = {fmt0_recB_rawIn_sign,_fmt0_recB_T_4,fmt0_recB_rawIn__sExp[20:0]}; // @[recFNFromFN.scala 49:45]
  wire  divOutValid = divsqrt_f0_io_outValid_div; // @[Emitscientist.scala 47:48]
  reg  busy; // @[Emitscientist.scala 52:21]
  wire  _T = ~io_opSel; // @[Emitscientist.scala 54:20]
  reg  divPending; // @[Emitscientist.scala 56:33]
  wire  _GEN_0 = ~busy & _T | divPending; // @[Emitscientist.scala 57:43 58:22 56:33]
  wire  _GEN_2 = divPending & divsqrt_f0_io_inReady | busy; // @[Emitscientist.scala 61:51 63:16 52:21]
  wire [512:0] outRec = ~io_opSel ? divsqrt_f0_io_out : 513'h0; // @[Emitscientist.scala 54:20 65:16 48:27]
  wire  recNonZero = |outRec; // @[Emitscientist.scala 72:27]
  wire [23:0] outIeee_rawIn_exp = outRec[511:488]; // @[rawFloatFromRecFN.scala 51:21]
  wire  outIeee_rawIn_isZero = outIeee_rawIn_exp[23:21] == 3'h0; // @[rawFloatFromRecFN.scala 52:53]
  wire  outIeee_rawIn_isSpecial = outIeee_rawIn_exp[23:22] == 2'h3; // @[rawFloatFromRecFN.scala 53:53]
  wire  outIeee_rawIn__isNaN = outIeee_rawIn_isSpecial & outIeee_rawIn_exp[21]; // @[rawFloatFromRecFN.scala 56:33]
  wire  outIeee_rawIn__isInf = outIeee_rawIn_isSpecial & ~outIeee_rawIn_exp[21]; // @[rawFloatFromRecFN.scala 57:33]
  wire  outIeee_rawIn__sign = outRec[512]; // @[rawFloatFromRecFN.scala 59:25]
  wire [24:0] outIeee_rawIn__sExp = {1'b0,$signed(outIeee_rawIn_exp)}; // @[rawFloatFromRecFN.scala 60:27]
  wire  _outIeee_rawIn_out_sig_T = ~outIeee_rawIn_isZero; // @[rawFloatFromRecFN.scala 61:35]
  wire [489:0] outIeee_rawIn__sig = {1'h0,_outIeee_rawIn_out_sig_T,outRec[487:0]}; // @[rawFloatFromRecFN.scala 61:44]
  wire  outIeee_isSubnormal = $signed(outIeee_rawIn__sExp) < 25'sh400002; // @[fNFromRecFN.scala 51:38]
  wire [8:0] outIeee_denormShiftDist = 9'h1 - outIeee_rawIn__sExp[8:0]; // @[fNFromRecFN.scala 52:35]
  wire [488:0] _outIeee_denormFract_T_1 = outIeee_rawIn__sig[489:1] >> outIeee_denormShiftDist; // @[fNFromRecFN.scala 53:42]
  wire [487:0] outIeee_denormFract = _outIeee_denormFract_T_1[487:0]; // @[fNFromRecFN.scala 53:60]
  wire [22:0] _outIeee_expOut_T_2 = outIeee_rawIn__sExp[22:0] - 23'h400001; // @[fNFromRecFN.scala 58:45]
  wire [22:0] _outIeee_expOut_T_3 = outIeee_isSubnormal ? 23'h0 : _outIeee_expOut_T_2; // @[fNFromRecFN.scala 56:16]
  wire  _outIeee_expOut_T_4 = outIeee_rawIn__isNaN | outIeee_rawIn__isInf; // @[fNFromRecFN.scala 60:44]
  wire [22:0] _outIeee_expOut_T_6 = _outIeee_expOut_T_4 ? 23'h7fffff : 23'h0; // @[Bitwise.scala 77:12]
  wire [22:0] outIeee_expOut = _outIeee_expOut_T_3 | _outIeee_expOut_T_6; // @[fNFromRecFN.scala 60:15]
  wire [487:0] _outIeee_fractOut_T_1 = outIeee_rawIn__isInf ? 488'h0 : outIeee_rawIn__sig[487:0]; // @[fNFromRecFN.scala 64:20]
  wire [487:0] outIeee_fractOut = outIeee_isSubnormal ? outIeee_denormFract : _outIeee_fractOut_T_1; // @[fNFromRecFN.scala 62:16]
  wire [511:0] outIeee = {outIeee_rawIn__sign,outIeee_expOut,outIeee_fractOut}; // @[Cat.scala 33:92]
  DivSqrtRecFM_small_e23_s489 divsqrt_f0 ( // @[Emitscientist.scala 39:26]
    .clock(divsqrt_f0_clock),
    .reset(divsqrt_f0_reset),
    .io_inReady(divsqrt_f0_io_inReady),
    .io_inValid(divsqrt_f0_io_inValid),
    .io_a(divsqrt_f0_io_a),
    .io_b(divsqrt_f0_io_b),
    .io_roundingMode(divsqrt_f0_io_roundingMode),
    .io_outValid_div(divsqrt_f0_io_outValid_div),
    .io_out(divsqrt_f0_io_out),
    .io_exceptionFlags(divsqrt_f0_io_exceptionFlags)
  );
  assign io_out = recNonZero ? outIeee : 512'h0; // @[Emitscientist.scala 75:16]
  assign io_exceptionFlags = ~io_opSel ? divsqrt_f0_io_exceptionFlags : 5'h0; // @[Emitscientist.scala 54:20 66:16 50:27]
  assign divsqrt_f0_clock = clock;
  assign divsqrt_f0_reset = reset;
  assign divsqrt_f0_io_inValid = ~io_opSel & divPending; // @[Emitscientist.scala 54:20 60:19 40:27]
  assign divsqrt_f0_io_a = {_fmt0_recA_T_7,fmt0_recA_rawIn__sig[487:0]}; // @[recFNFromFN.scala 50:41]
  assign divsqrt_f0_io_b = {_fmt0_recB_T_7,fmt0_recB_rawIn__sig[487:0]}; // @[recFNFromFN.scala 50:41]
  assign divsqrt_f0_io_roundingMode = roundingMatches_0 ? io_roundingMode : 3'h0; // @[Emitscientist.scala 21:25]
  always @(posedge clock) begin
    if (reset) begin // @[Emitscientist.scala 52:21]
      busy <= 1'h0; // @[Emitscientist.scala 52:21]
    end else if (~io_opSel) begin // @[Emitscientist.scala 54:20]
      if (divOutValid) begin // @[Emitscientist.scala 68:27]
        busy <= 1'h0; // @[Emitscientist.scala 68:34]
      end else begin
        busy <= _GEN_2;
      end
    end
    if (reset) begin // @[Emitscientist.scala 56:33]
      divPending <= 1'h0; // @[Emitscientist.scala 56:33]
    end else if (divPending & divsqrt_f0_io_inReady) begin // @[Emitscientist.scala 61:51]
      divPending <= 1'h0; // @[Emitscientist.scala 62:22]
    end else begin
      divPending <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  divPending = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
